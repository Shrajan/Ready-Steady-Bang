////////////////////////////////////////////////////////////////////////////////
 /*
 FPGA Project Name     : Ready Steady Bang
 Top level Entity Name : Video_Engine
 Target Device		   : Cyclone V
 
 Code Authors          : Sanjith Chandran and Shrajan Bhandary 
 Date Created          : 20/04/2019 
 Location 			   : University of Leeds
 Module 			   : ELEC5566M FPGA Design for System-on-chip
 
 -------------------------------------------------------------------------------
 
 Description of the Verilog Module: 
	The module defines the values of pixels for different states of the game.
 
 */
//////////////////////////////////////////////////////////////////////////////// 

/* ceil(log2(N)) Preprocessor Macro */
`define clog2(x) ( \
	((x) <= 2) ? 1 : \
	((x) <= 4) ? 2 : \
	((x) <= 8) ? 3 : \
	((x) <= 16) ? 4 : \
	((x) <= 32) ? 5 : \
	((x) <= 64) ? 6 : \
	((x) <= 128) ? 7 : \
	((x) <= 256) ? 8 : \
	((x) <= 512) ? 9 : \
	((x) <= 1024) ? 10 : \
	((x) <= 2048) ? 11 : \
	((x) <= 4096) ? 12 : 16)

module Video_Engine #(															// Start of the module.

    /* Parameter List of the Video_Engine */
    parameter LCD_WIDTH  	      = 240				      ,						// The number of pixels in the x-direction is 240.
	parameter LCD_HEIGHT 	      = 320				      ,						// The number of pixels in the y-direction is 320.
	parameter X_ADDRESS_WIDTH     = `clog2(LCD_WIDTH)     ,						// Number of bits required to store the x-address.
	parameter Y_ADDRESS_WIDTH 	  = `clog2(LCD_HEIGHT)    ,						// Number of bits required to store the y-address.
	
	parameter NO_GAME_STATES	  = 35				      ,						// The number of possible states (Screens).
	parameter STATE_ADDRESS_WIDTH = `clog2(NO_GAME_STATES),						// Number of bits required to store the different number of states.
	
	parameter PIXEL_ADDRESS_WIDTH = 16                    ,						// Number of bits required to colour a pixel.
	parameter PLAYER_ID			  = 1											// The ID is either 1 or 2 depending on the board that the program runs.
)(
	/* Port List of the Video_Engine */
    input 	  [(X_ADDRESS_WIDTH-1):0] lcd_pixel_x_address	,					// The current x-coordinate of the LCD pixel.	
	input 	  [(Y_ADDRESS_WIDTH-1):0] lcd_pixel_y_address	,					// The current y-coordinate of the LCD pixel.
	input 	  [(STATE_ADDRESS_WIDTH-1):0] game_states     	,					// The current state of the game screen.
	output 	  reg [(PIXEL_ADDRESS_WIDTH-1):0] lcd_pixel_data					// The data values that determine the colour of the pixel.
);	
	/* Local Parameters list containing the screen states of LCD of the Game_Engine.*/
	/* States that determine the settings of the game.*/
	localparam A_STATE = 6'b000001;												// Main screen of the game.
	localparam B_STATE = 6'b000010;												// One player version screen of the game.
	localparam C_STATE = 6'b000011;												// Two player version screen of the game.
	
	/* States that control one player version of the game.*/
	localparam D_1_STATE = 6'b000100;											// Start screen of the One player version of the game.
	localparam E_1_STATE = 6'b000101;											// Empty screen 1 of the One player version of the game.
	localparam F_1_STATE = 6'b000110;											// Ready screen of the One player version of the game.
	localparam G_1_STATE = 6'b000111;											// Empty screen 2 of the One player version of the game.
	localparam H_1_STATE = 6'b001000;											// Steady screen of the One player version of the game.
	localparam I_1_STATE = 6'b001001;											// Empty screen 3 of the One player version of the game.
	localparam J_1_STATE = 6'b001010;											// Bang screen of the One player version of the game.
	localparam K_1_STATE = 6'b001011;											// First Player kill screen of the One player version of the game.
	localparam L_1_STATE = 6'b001100;											// Second Player kill screen of the One player version of the game.
	localparam M_1_STATE = 6'b001101;											// Both Player kill screen of the One player version of the game.
	localparam N_1_STATE = 6'b001110;											// Next - First Player kill screen of the One player version of the game.
	localparam O_1_STATE = 6'b001111;											// Next - Second Player kill screen of the One player version of the game.
	localparam P_1_STATE = 6'b010000;											// Next - Both Player kill screen of the One player version of the game.
	localparam Q_1_STATE = 6'b010001;											// Player one Winner screen of the One player version of the game.
	localparam R_1_STATE = 6'b010010;											// Player two Winner screen of the One player version of the game.
	
	/* States that control two player version of the game.*/
	localparam D_2_STATE = 6'b010100;											// Start screen of the Two player version of the game.
	localparam E_2_STATE = 6'b010101;											// Empty screen 1 of the Two player version of the game.
	localparam F_2_STATE = 6'b010110;											// Ready screen of the Two player version of the game.
	localparam G_2_STATE = 6'b010111;											// Empty screen 2 of the Two player version of the game.
	localparam H_2_STATE = 6'b011000;											// Steady screen of the Two player version of the game.
	localparam I_2_STATE = 6'b011001;											// Empty screen 3 of the Two player version of the game.
	localparam J_2_STATE = 6'b011010;											// Bang screen of the Two player version of the game.
	localparam K_2_STATE = 6'b011011;											// First Player kill screen of the Two player version of the game.
	localparam L_2_STATE = 6'b011100;											// Second Player kill screen of the Two player version of the game.
	localparam M_2_STATE = 6'b011101;											// Both Player kill screen of the Two player version of the game.
	localparam N_2_STATE = 6'b011110;											// Next - First Player kill screen of the Two player version of the game.
	localparam O_2_STATE = 6'b011111;											// Next - Second Player kill screen of the Two player version of the game.
	localparam P_2_STATE = 6'b100000;											// Next - Both Player kill screen of the Two player version of the game.
	localparam Q_2_STATE = 6'b100001;											// Player one Winner screen of the Two player version of the game.
	localparam R_2_STATE = 6'b100010;											// Player two Winner screen of the Two player version of the game.
	
	always @ ( game_states, lcd_pixel_y_address, lcd_pixel_x_address )
		begin 
		
			if ( PLAYER_ID == 1 )
				begin
					localparam SCARF_COLOUR = 16'h07E0;
					localparam SCARF2_COLOUR = 16'hF81F;
					
					/* Beginning of Main screen of the game. */
					if ( game_states == A_STATE  )
						begin
						
							localparam READY_X = 100;
							localparam READY_Y = 130;
							localparam READY_COLOUR = 16'hFFFF;
							localparam STEADY_X = 95;
							localparam STEADY_Y = 150;
							localparam STEADY_COLOUR = 16'hFFFF;
							localparam BANG_X = 105;
							localparam BANG_Y = 170;
							localparam BANG_COLOUR = 16'hFFFF;

							//1P
							localparam GUNMAN_X = 85;
							localparam GUNMAN_Y = 200;
							localparam BODY_COLOUR = 16'hFFFF;
							localparam BOX_COLOUR = 16'hFFFF;
							////localparam SCARF_COLOUR = 16'h07E0;
							localparam BELT_COLOUR = 16'hDA22;
							localparam GUN_COLOUR = 16'hA516;
							localparam PANTS_COLOUR = 16'h001F;
							localparam EXPLODE = 16'hF800;

							//2P
							localparam GUNMAN2_X = 145;
							localparam GUNMAN2_Y = 200;
							localparam BODY2_COLOUR = 16'hFFFF;
							localparam BOX2_COLOUR = 16'hFFFF;
							//localparam SCARF2_COLOUR = 16'hF81F;
							localparam BELT2_COLOUR = 16'hDA22;
							localparam GUN2_COLOUR = 16'hA516;
							localparam PANTS2_COLOUR = 16'h001F;
							localparam EXPLODE2 = 16'hF800;
							
							//WORD READY
							//READY=30
							
							//Letter R
							if (((lcd_pixel_y_address >= READY_Y) && (lcd_pixel_y_address <= (READY_Y+15)))&& (lcd_pixel_x_address == READY_X))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
								
							else if (((lcd_pixel_x_address >=READY_X) && (lcd_pixel_x_address <= (READY_X+7)))&& (lcd_pixel_y_address == READY_Y))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= (READY_Y+7)))&& (lcd_pixel_x_address == (READY_X+7)))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >= READY_X) && (lcd_pixel_x_address <= (READY_X+7)))&& (lcd_pixel_y_address == (READY_Y+7)))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if ((lcd_pixel_x_address==READY_X+1) && (lcd_pixel_y_address==READY_Y+9))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==READY_X+2) && (lcd_pixel_y_address==READY_Y+10))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==READY_X+3) && (lcd_pixel_y_address==READY_Y+11)) 
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==READY_X+4) && (lcd_pixel_y_address==READY_Y+12))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==READY_X+5) && (lcd_pixel_y_address==READY_Y+13))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==READY_X+6) && (lcd_pixel_y_address==READY_Y+14))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==READY_X+7) && (lcd_pixel_y_address==READY_Y+15))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	 
								end
								
							//Letter E
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+10))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y+7))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y+15))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
								
							//Letter A
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+20))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=READY_X+20) && (lcd_pixel_x_address <= READY_X+27))&& (lcd_pixel_y_address == READY_Y))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+20) && (lcd_pixel_x_address <= READY_X+27))&& (lcd_pixel_y_address == READY_Y+7))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+27))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
								
							//Letter D
							else if (((lcd_pixel_y_address >=READY_Y+4) && (lcd_pixel_y_address <= READY_Y+11))&& (lcd_pixel_x_address == READY_X+37))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+30))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+30) && (lcd_pixel_x_address <= READY_X+33))&& (lcd_pixel_y_address == READY_Y))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+30) && (lcd_pixel_x_address <= READY_X+33))&& (lcd_pixel_y_address == READY_Y+15))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if ((lcd_pixel_x_address==READY_X+33)  && (lcd_pixel_y_address==READY_Y))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if ((lcd_pixel_x_address==READY_X+33)  && (lcd_pixel_y_address==READY_Y+15))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if ((lcd_pixel_x_address==READY_X+34) && (lcd_pixel_y_address==READY_Y+1))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==READY_X+34) && (lcd_pixel_y_address==READY_Y+14))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==READY_X+35) && (lcd_pixel_y_address==READY_Y+2))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if ((lcd_pixel_x_address==READY_X+35) && (lcd_pixel_y_address==READY_Y+13))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if ((lcd_pixel_x_address==READY_X+36) && (lcd_pixel_y_address==READY_Y+3))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if ((lcd_pixel_x_address==READY_X+36) && (lcd_pixel_y_address==READY_Y+12))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							
							//Letter Y
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+47))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+7))&& (lcd_pixel_x_address == READY_X+40))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
								
							else if (((lcd_pixel_x_address >=READY_X+40) && (lcd_pixel_x_address <= READY_X+47))&& (lcd_pixel_y_address == READY_Y+7))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+40) && (lcd_pixel_x_address <= READY_X+47))&& (lcd_pixel_y_address == READY_Y+15))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							
							
							//STEADY_Y+ & STEADY_X+
							//STEADY_COLOUR
							//Letter S
							//else
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+7))&& (lcd_pixel_x_address == STEADY_X))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y+7))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y+15))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=STEADY_Y+8) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+7))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
								
								//Letter T
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+14))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STEADY_X+10) && (lcd_pixel_x_address <= STEADY_X+17))&& (lcd_pixel_y_address == STEADY_Y))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							
							//Letter E
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+20))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y+7))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y+15))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							
							//Letter A
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+30))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STEADY_X+30) && (lcd_pixel_x_address <= STEADY_X+37))&& (lcd_pixel_y_address == STEADY_Y))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+30) && (lcd_pixel_x_address <= STEADY_X+37))&& (lcd_pixel_y_address == STEADY_Y+7))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+37))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
								
							//Letter D
							else if (((lcd_pixel_y_address >=STEADY_Y+4) && (lcd_pixel_y_address <= STEADY_Y+11))&& (lcd_pixel_x_address == STEADY_X+47))
								begin
									lcd_pixel_data[15:0] <=STEADY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+40))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+40) && (lcd_pixel_x_address <= STEADY_X+43))&& (lcd_pixel_y_address == STEADY_Y))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+40) && (lcd_pixel_x_address <= STEADY_X+43))&& (lcd_pixel_y_address == STEADY_Y+15))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+43) && (lcd_pixel_y_address == STEADY_Y))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==STEADY_X+43) && (lcd_pixel_y_address == STEADY_Y+15))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==STEADY_X+44) && (lcd_pixel_y_address == STEADY_Y+1))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+44) && (lcd_pixel_y_address == STEADY_Y+14))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+45) && (lcd_pixel_y_address == STEADY_Y+2))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+45) && (lcd_pixel_y_address == STEADY_Y+13))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+46) && (lcd_pixel_y_address == STEADY_Y+3))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+46) && (lcd_pixel_y_address == STEADY_Y+12))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							
							//Letter Y
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+57))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+7))&& (lcd_pixel_x_address == STEADY_X+50))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
								
							else if (((lcd_pixel_x_address >=STEADY_X+50) && (lcd_pixel_x_address <= STEADY_X+57))&& (lcd_pixel_y_address == STEADY_Y+7))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+50) && (lcd_pixel_x_address <= STEADY_X+57))&& (lcd_pixel_y_address == STEADY_Y+15))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
								
							
							//BANG_Y+=70
							//BANG_X+=30
							//BANG_COLOUR
							//Letter B
							else if (((lcd_pixel_y_address >=BANG_Y+3) && (lcd_pixel_y_address <= BANG_Y+4))&& (lcd_pixel_x_address == BANG_X+7))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_y_address >=BANG_Y+10) && (lcd_pixel_y_address <= BANG_Y+12))&& (lcd_pixel_x_address == BANG_X+7))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
								
							else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y+7))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y+15))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+1))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+6))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+8))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+14))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
								
							else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+2))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+5))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+9))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+13))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							//Letter A
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+10))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=BANG_X+10) && (lcd_pixel_x_address <= BANG_X+17))&& (lcd_pixel_y_address == BANG_Y))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_x_address >=BANG_X+10) && (lcd_pixel_x_address <= BANG_X+17))&& (lcd_pixel_y_address == BANG_Y+7))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+17))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
								
							//Letter N
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+20))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+27))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+1))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+2))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+3))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+3))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+4))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+5))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+5))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+6))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+7))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end

							
							else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+7))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+8))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+9))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+9))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+10))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+11))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							
							
							else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+11))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+12))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+13))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							
							//Letter G
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+30))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=BANG_X+30) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_x_address >=BANG_X+34) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y+7))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_x_address >=BANG_X+30) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y+15))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_y_address >=BANG_Y+7) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+37))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end						
							
							//HEAD
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							
							//Gunman Body
							
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end	
								
							//HEAD
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							
							//GUNMAN2 Body
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end	
							else 	
								begin
									lcd_pixel_data <= 16'h0000;
								end
							
						end 
						/* End of Main screen of the game. */
					
					/*Selecting 1-Player Mode*/
					else if ( game_states == B_STATE )
						begin
						
						localparam LCD_WIDTH  = 240;
						localparam LCD_HEIGHT = 320;

						//1P
						localparam GUNMAN_X = 50;
						localparam GUNMAN_Y = 150;
						localparam BODY_COLOUR = 16'h0000;
						//localparam SCARF_COLOUR = 16'h07E0;
						localparam BELT_COLOUR = 16'hDA22;
						localparam GUN_COLOUR = 16'hA516;
						localparam PANTS_COLOUR = 16'h001F;
						localparam EXPLODE = 16'hF800;

						//2P
						localparam GUNMAN2_X = 130;
						localparam GUNMAN2_Y = 150;
						localparam BODY2_COLOUR = 16'h0000;
						//localparam SCARF2_COLOUR = 16'hF81F;
						localparam BELT2_COLOUR = 16'hDA22;
						localparam GUN2_COLOUR = 16'hA516;
						localparam PANTS2_COLOUR = 16'h001F;
						localparam EXPLODE2 = 16'hF800;


						localparam _1P_X = 53;
						localparam _1P_Y = 120;
						localparam _1P_COLOUR = 16'h0000;

						localparam _2P_X = 150;
						localparam _2P_Y = 120;
						localparam _2P_COLOUR = 16'h0000;

						localparam BOX_COLOUR = 16'h0000;
						localparam BOX2_COLOUR = 16'h0000;


								//Player One
									//1
								if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+1))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+2))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+3))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if ((lcd_pixel_x_address==_1P_X+3) && (lcd_pixel_y_address == _1P_Y))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+3) && (lcd_pixel_y_address == _1P_Y+1))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+3))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+4))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+5))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
									
								else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= _1P_Y+15))&& (lcd_pixel_x_address == _1P_X+4))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >=_1P_X) && (lcd_pixel_x_address <= _1P_X+8))&& (lcd_pixel_y_address == _1P_Y+15))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								//P	
								else if (((lcd_pixel_y_address >= _1P_Y) && (lcd_pixel_y_address <= (_1P_Y+15)))&& (lcd_pixel_x_address == _1P_X+10))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if (((lcd_pixel_x_address >=_1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == _1P_Y))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= (_1P_Y+7)))&& (lcd_pixel_x_address == (_1P_X+17)))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >= _1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == (_1P_Y+7)))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
									
								//PLAYER 2
							
								else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= _2P_Y+7))&& (lcd_pixel_x_address == _2P_X+7))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y+7))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y+15))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_y_address >=_2P_Y+8) && (lcd_pixel_y_address <= _2P_Y+15))&& (lcd_pixel_x_address == _2P_X))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_y_address >= _2P_Y) && (lcd_pixel_y_address <= (_2P_Y+15)))&& (lcd_pixel_x_address == _2P_X+10))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
									
								else if (((lcd_pixel_x_address >=_2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == _2P_Y))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= (_2P_Y+7)))&& (lcd_pixel_x_address == (_2P_X+17)))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >= _2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == (_2P_Y+7)))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								//
								//
								
								//Gunman 1
								
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end

								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT_COLOUR;
									end
								
								//Gunman Body
								
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end	
								
								//BOX for P1
								else if (((lcd_pixel_y_address >=(GUNMAN_Y-5)) && (lcd_pixel_y_address <= (GUNMAN_Y+38)))&&(lcd_pixel_x_address == (GUNMAN_X-8)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end	
								else if (((lcd_pixel_y_address >=(GUNMAN_Y-5)) && (lcd_pixel_y_address <= (GUNMAN_Y+38)))&&(lcd_pixel_x_address == (GUNMAN_X+26)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X-8) && (lcd_pixel_x_address <= (GUNMAN_X+26)))&&(lcd_pixel_y_address == (GUNMAN_Y-5)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X-8) && (lcd_pixel_x_address <= (GUNMAN_X+26)))&&(lcd_pixel_y_address == (GUNMAN_Y+38)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end	
									
								//2P 
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
							
								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								
								//GUNMAN2 Body
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end	
									
								//DUPLICATE FOR SELECTING OPTION	
										
								
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+47)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+50)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+47)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+50)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+45)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+52)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+45)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+52)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+48)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+49)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+46) && (lcd_pixel_x_address <= (GUNMAN2_X+51)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+46) && (lcd_pixel_x_address <= (GUNMAN2_X+51)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+48) && (lcd_pixel_x_address <= (GUNMAN2_X+49)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+48) && (lcd_pixel_x_address <= (GUNMAN2_X+49)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								
								//GUNMAN2 Body
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN2_X+39) && (lcd_pixel_x_address >= (GUNMAN2_X+38)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN2_X+39) && (lcd_pixel_x_address >= (GUNMAN2_X+38)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+58) && (lcd_pixel_x_address <= (GUNMAN2_X+59)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+58) && (lcd_pixel_x_address <= (GUNMAN2_X+59)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+37)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+36)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+60)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+61)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+40)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+41)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+42)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+43)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+56)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+57)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+54)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+44)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+45)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+52)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+53)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+42)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+43)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+41)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+54)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end	

								else 	
									begin
										//lcd_pixel_data <= 16'hFFFF;
										lcd_pixel_data <= 16'hFFFF;
									end

						end
					/*End of Selecting 1-Player Mode*/
					
					/*Selecting 2-Player Mode*/
					else if ( game_states == C_STATE )
						begin
											
						localparam LCD_WIDTH  = 240;
						localparam LCD_HEIGHT = 320;

						//1P
						localparam GUNMAN_X = 50;
						localparam GUNMAN_Y = 150;
						localparam BODY_COLOUR = 16'h0000;
						//localparam SCARF_COLOUR = 16'h07E0;
						localparam BELT_COLOUR = 16'hDA22;
						localparam GUN_COLOUR = 16'hA516;
						localparam PANTS_COLOUR = 16'h001F;
						localparam EXPLODE = 16'hF800;

						//2P
						localparam GUNMAN2_X = 130;
						localparam GUNMAN2_Y = 150;
						localparam BODY2_COLOUR = 16'h0000;
						//localparam SCARF2_COLOUR = 16'hF81F;
						localparam BELT2_COLOUR = 16'hDA22;
						localparam GUN2_COLOUR = 16'hA516;
						localparam PANTS2_COLOUR = 16'h001F;
						localparam EXPLODE2 = 16'hF800;


						localparam _1P_X = 53;
						localparam _1P_Y = 120;
						localparam _1P_COLOUR = 16'h0000;

						localparam _2P_X = 150;
						localparam _2P_Y = 120;
						localparam _2P_COLOUR = 16'h0000;

						localparam BOX_COLOUR = 16'h0000;
						localparam BOX2_COLOUR = 16'h0000;



								if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+1))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+2))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+3))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if ((lcd_pixel_x_address==_1P_X+3) && (lcd_pixel_y_address == _1P_Y))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+3) && (lcd_pixel_y_address == _1P_Y+1))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+3))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+4))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+5))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
									
								else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= _1P_Y+15))&& (lcd_pixel_x_address == _1P_X+4))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >=_1P_X) && (lcd_pixel_x_address <= _1P_X+8))&& (lcd_pixel_y_address == _1P_Y+15))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								//P	
								else if (((lcd_pixel_y_address >= _1P_Y) && (lcd_pixel_y_address <= (_1P_Y+15)))&& (lcd_pixel_x_address == _1P_X+10))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if (((lcd_pixel_x_address >=_1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == _1P_Y))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= (_1P_Y+7)))&& (lcd_pixel_x_address == (_1P_X+17)))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >= _1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == (_1P_Y+7)))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
									
								//PLAYER 2
							
								else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= _2P_Y+7))&& (lcd_pixel_x_address == _2P_X+7))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y+7))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y+15))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_y_address >=_2P_Y+8) && (lcd_pixel_y_address <= _2P_Y+15))&& (lcd_pixel_x_address == _2P_X))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_y_address >= _2P_Y) && (lcd_pixel_y_address <= (_2P_Y+15)))&& (lcd_pixel_x_address == _2P_X+10))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
									
								else if (((lcd_pixel_x_address >=_2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == _2P_Y))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= (_2P_Y+7)))&& (lcd_pixel_x_address == (_2P_X+17)))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >= _2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == (_2P_Y+7)))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								//
								//
								
								//Gunman 1
								
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end

								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT_COLOUR;
									end
								
								//Gunman Body
								
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end	
								
								/*//BOX for P1
								else if (((lcd_pixel_y_address >=(GUNMAN_Y-5)) && (lcd_pixel_y_address <= (GUNMAN_Y+38)))&&(lcd_pixel_x_address == (GUNMAN_X-8)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end	
								else if (((lcd_pixel_y_address >=(GUNMAN_Y-5)) && (lcd_pixel_y_address <= (GUNMAN_Y+38)))&&(lcd_pixel_x_address == (GUNMAN_X+26)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X-8) && (lcd_pixel_x_address <= (GUNMAN_X+26)))&&(lcd_pixel_y_address == (GUNMAN_Y-5)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X-8) && (lcd_pixel_x_address <= (GUNMAN_X+26)))&&(lcd_pixel_y_address == (GUNMAN_Y+38)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end*/	
									
								//2P 
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
							
								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								
								//GUNMAN2 Body
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end	
									
								//DUPLICATE FOR SELECTING OPTION	
										
								
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+47)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+50)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+47)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+50)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+45)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+52)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+45)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+52)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+48)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+49)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+46) && (lcd_pixel_x_address <= (GUNMAN2_X+51)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+46) && (lcd_pixel_x_address <= (GUNMAN2_X+51)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+48) && (lcd_pixel_x_address <= (GUNMAN2_X+49)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+48) && (lcd_pixel_x_address <= (GUNMAN2_X+49)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								
								//GUNMAN2 Body
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN2_X+39) && (lcd_pixel_x_address >= (GUNMAN2_X+38)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN2_X+39) && (lcd_pixel_x_address >= (GUNMAN2_X+38)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+58) && (lcd_pixel_x_address <= (GUNMAN2_X+59)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+58) && (lcd_pixel_x_address <= (GUNMAN2_X+59)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+37)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+36)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+60)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+61)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+40)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+41)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+42)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+43)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+56)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+57)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+54)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+44)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+45)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+52)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+53)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+42)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+43)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+41)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+54)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end	
								
								//BOX for P2
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y-5)) && (lcd_pixel_y_address <= (GUNMAN2_Y+38)))&&(lcd_pixel_x_address == (GUNMAN2_X-8)))
									begin
										lcd_pixel_data[15:0] <= BOX2_COLOUR;
									end	
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y-5)) && (lcd_pixel_y_address <= (GUNMAN2_Y+38)))&&(lcd_pixel_x_address == (GUNMAN2_X+66)))
									begin
										lcd_pixel_data[15:0] <= BOX2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X-8) && (lcd_pixel_x_address <= (GUNMAN2_X+66)))&&(lcd_pixel_y_address == (GUNMAN2_Y-5)))
									begin
										lcd_pixel_data[15:0] <= BOX2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X-8) && (lcd_pixel_x_address <= (GUNMAN2_X+66)))&&(lcd_pixel_y_address == (GUNMAN2_Y+38)))
									begin
										lcd_pixel_data[15:0] <= BOX2_COLOUR;
									end
									
								
								else 	
									begin
										//lcd_pixel_data <= 16'hFFFF;
										lcd_pixel_data <= 16'hFFFF;
									end
								  
							
											
									
						end
					/*End of Selecting 2-Player Mode*/
					
					/* Beginning of Select Player screen. */
					else if ( game_states == D_1_STATE || game_states == D_2_STATE  )
						begin
						
							localparam LCD_WIDTH  = 240;
							localparam LCD_HEIGHT = 320;

							localparam STARTGAME_X = 105;
							localparam STARTGAME_Y = 150;
							localparam STARTGAME_COLOUR = 16'h0000;

							//1P
							localparam GUNMAN_X = 115;
							localparam GUNMAN_Y = 250;
							localparam BODY_COLOUR = 16'h0000;
							//localparam SCARF_COLOUR = 16'h07E0;
							localparam BELT_COLOUR = 16'hDA22;
							localparam GUN_COLOUR = 16'hA516;
							localparam PANTS_COLOUR = 16'h001F;
							localparam EXPLODE = 16'hF800;

							//2P
							localparam GUNMAN2_X = 115;
							localparam GUNMAN2_Y = 50;
							localparam BODY2_COLOUR = 16'h0000;
							//localparam SCARF2_COLOUR = 16'hF81F;
							localparam BELT2_COLOUR = 16'hDA22;
							localparam GUN2_COLOUR = 16'hA516;
							localparam PANTS2_COLOUR = 16'h001F;
							localparam EXPLODE2 = 16'hF800;
							
							//STARTGAME_Y+ & STARTGAME_X+
							//STARTGAME_COLOUR
							//Letter S
							//else
							if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= STARTGAME_Y+7))&& (lcd_pixel_x_address == STARTGAME_X))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STARTGAME_X) && (lcd_pixel_x_address <= STARTGAME_X+7))&& (lcd_pixel_y_address == STARTGAME_Y))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STARTGAME_X) && (lcd_pixel_x_address <= STARTGAME_X+7))&& (lcd_pixel_y_address == STARTGAME_Y+7))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STARTGAME_X) && (lcd_pixel_x_address <= STARTGAME_X+7))&& (lcd_pixel_y_address == STARTGAME_Y+15))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if (((lcd_pixel_y_address >=STARTGAME_Y+8) && (lcd_pixel_y_address <= STARTGAME_Y+15))&& (lcd_pixel_x_address == STARTGAME_X+7))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
								
								//Letter T
							else if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= STARTGAME_Y+15))&& (lcd_pixel_x_address == STARTGAME_X+14))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STARTGAME_X+10) && (lcd_pixel_x_address <= STARTGAME_X+17))&& (lcd_pixel_y_address == STARTGAME_Y))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							
							
							//Letter A
							else if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= STARTGAME_Y+15))&& (lcd_pixel_x_address == STARTGAME_X+20))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STARTGAME_X+20) && (lcd_pixel_x_address <= STARTGAME_X+27))&& (lcd_pixel_y_address == STARTGAME_Y))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STARTGAME_X+20) && (lcd_pixel_x_address <= STARTGAME_X+27))&& (lcd_pixel_y_address == STARTGAME_Y+7))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= STARTGAME_Y+15))&& (lcd_pixel_x_address == STARTGAME_X+27))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
								
							//Letter R
							else if (((lcd_pixel_y_address >= STARTGAME_Y) && (lcd_pixel_y_address <= (STARTGAME_Y+15)))&& (lcd_pixel_x_address == STARTGAME_X+30))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
								
							else if (((lcd_pixel_x_address >=STARTGAME_X+30) && (lcd_pixel_x_address <= (STARTGAME_X+37)))&& (lcd_pixel_y_address == STARTGAME_Y))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= (STARTGAME_Y+7)))&& (lcd_pixel_x_address == (STARTGAME_X+37)))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end	
							else if (((lcd_pixel_x_address >= STARTGAME_X+30) && (lcd_pixel_x_address <= (STARTGAME_X+37)))&& (lcd_pixel_y_address == (STARTGAME_Y+7)))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+31) && (lcd_pixel_y_address==STARTGAME_Y+9))
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+32) && (lcd_pixel_y_address==STARTGAME_Y+10))
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+33) && (lcd_pixel_y_address==STARTGAME_Y+11)) 
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+34) && (lcd_pixel_y_address==STARTGAME_Y+12))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+35) && (lcd_pixel_y_address==STARTGAME_Y+13))
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+36) && (lcd_pixel_y_address==STARTGAME_Y+14))
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+37) && (lcd_pixel_y_address==STARTGAME_Y+15))
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	 
								end
							//Letter T
							else if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= STARTGAME_Y+15))&& (lcd_pixel_x_address == STARTGAME_X+44))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STARTGAME_X+40) && (lcd_pixel_x_address <= STARTGAME_X+47))&& (lcd_pixel_y_address == STARTGAME_Y))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							
							
							//HEAD
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end

							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							
							//Gunman Body
							
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end	
							
								
								
							
							//HEAD
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//scarf 
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							
							//GUNMAN2 Body
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end	
							else 	
								begin	
									lcd_pixel_data <= 16'hFFFF;
								end
							
						end 
						/* End of Select Player screen. */
					
					/*In-Between Screens*/
					else if ( game_states == E_1_STATE || game_states == G_1_STATE || game_states == I_1_STATE || game_states == E_2_STATE || game_states == G_2_STATE || game_states == I_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				//HEAD
				if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
		   
						
						end
					/*End of In-Between Screens*/
					
					/*Ready Screen for Game*/
					else if ( game_states == F_1_STATE || game_states == F_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		localparam READY_X = 105;
		localparam READY_Y = 150;
		localparam READY_COLOUR = 16'h0000;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				//Letter R
				if (((lcd_pixel_y_address >= READY_Y) && (lcd_pixel_y_address <= (READY_Y+15)))&& (lcd_pixel_x_address == READY_X))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=READY_X) && (lcd_pixel_x_address <= (READY_X+7)))&& (lcd_pixel_y_address == READY_Y))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= (READY_Y+7)))&& (lcd_pixel_x_address == (READY_X+7)))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= READY_X) && (lcd_pixel_x_address <= (READY_X+7)))&& (lcd_pixel_y_address == (READY_Y+7)))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if ((lcd_pixel_x_address==READY_X+1) && (lcd_pixel_y_address==READY_Y+9))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==READY_X+2) && (lcd_pixel_y_address==READY_Y+10))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==READY_X+3) && (lcd_pixel_y_address==READY_Y+11)) 
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==READY_X+4) && (lcd_pixel_y_address==READY_Y+12))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==READY_X+5) && (lcd_pixel_y_address==READY_Y+13))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==READY_X+6) && (lcd_pixel_y_address==READY_Y+14))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==READY_X+7) && (lcd_pixel_y_address==READY_Y+15))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	 
					end
					
				//Letter E
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+10))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y+7))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y+15))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
					
				//Letter A
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+20))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=READY_X+20) && (lcd_pixel_x_address <= READY_X+27))&& (lcd_pixel_y_address == READY_Y))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+20) && (lcd_pixel_x_address <= READY_X+27))&& (lcd_pixel_y_address == READY_Y+7))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+27))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
					
				//Letter D
				else if (((lcd_pixel_y_address >=READY_Y+4) && (lcd_pixel_y_address <= READY_Y+11))&& (lcd_pixel_x_address == READY_X+37))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+30))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+30) && (lcd_pixel_x_address <= READY_X+33))&& (lcd_pixel_y_address == READY_Y))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+30) && (lcd_pixel_x_address <= READY_X+33))&& (lcd_pixel_y_address == READY_Y+15))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if ((lcd_pixel_x_address==READY_X+33)  && (lcd_pixel_y_address==READY_Y))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if ((lcd_pixel_x_address==READY_X+33)  && (lcd_pixel_y_address==READY_Y+15))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if ((lcd_pixel_x_address==READY_X+34) && (lcd_pixel_y_address==READY_Y+1))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==READY_X+34) && (lcd_pixel_y_address==READY_Y+14))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==READY_X+35) && (lcd_pixel_y_address==READY_Y+2))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if ((lcd_pixel_x_address==READY_X+35) && (lcd_pixel_y_address==READY_Y+13))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if ((lcd_pixel_x_address==READY_X+36) && (lcd_pixel_y_address==READY_Y+3))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if ((lcd_pixel_x_address==READY_X+36) && (lcd_pixel_y_address==READY_Y+12))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				
				//Letter Y
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+47))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+7))&& (lcd_pixel_x_address == READY_X+40))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=READY_X+40) && (lcd_pixel_x_address <= READY_X+47))&& (lcd_pixel_y_address == READY_Y+7))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+40) && (lcd_pixel_x_address <= READY_X+47))&& (lcd_pixel_y_address == READY_Y+15))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
			
						end
					/*End of Ready Screen for Game*/
					
					/*Steady Screen for Game*/
					else if (game_states == H_1_STATE || game_states == H_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		localparam STEADY_X = 105;
		localparam STEADY_Y = 150;
		localparam STEADY_COLOUR = 16'h0000;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+7))&& (lcd_pixel_x_address == STEADY_X))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y+7))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y+15))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=STEADY_Y+8) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+7))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
					
					//Letter T
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+14))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=STEADY_X+10) && (lcd_pixel_x_address <= STEADY_X+17))&& (lcd_pixel_y_address == STEADY_Y))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				
				//Letter E
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+20))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y+7))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y+15))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				
				//Letter A
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+30))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=STEADY_X+30) && (lcd_pixel_x_address <= STEADY_X+37))&& (lcd_pixel_y_address == STEADY_Y))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+30) && (lcd_pixel_x_address <= STEADY_X+37))&& (lcd_pixel_y_address == STEADY_Y+7))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+37))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
					
				//Letter D
				else if (((lcd_pixel_y_address >=STEADY_Y+4) && (lcd_pixel_y_address <= STEADY_Y+11))&& (lcd_pixel_x_address == STEADY_X+47))
					begin
						lcd_pixel_data[15:0] <=STEADY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+40))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+40) && (lcd_pixel_x_address <= STEADY_X+43))&& (lcd_pixel_y_address == STEADY_Y))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+40) && (lcd_pixel_x_address <= STEADY_X+43))&& (lcd_pixel_y_address == STEADY_Y+15))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+43) && (lcd_pixel_y_address == STEADY_Y))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==STEADY_X+43) && (lcd_pixel_y_address == STEADY_Y+15))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==STEADY_X+44) && (lcd_pixel_y_address == STEADY_Y+1))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+44) && (lcd_pixel_y_address == STEADY_Y+14))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+45) && (lcd_pixel_y_address == STEADY_Y+2))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+45) && (lcd_pixel_y_address == STEADY_Y+13))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+46) && (lcd_pixel_y_address == STEADY_Y+3))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+46) && (lcd_pixel_y_address == STEADY_Y+12))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				
				//Letter Y
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+57))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+7))&& (lcd_pixel_x_address == STEADY_X+50))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=STEADY_X+50) && (lcd_pixel_x_address <= STEADY_X+57))&& (lcd_pixel_y_address == STEADY_Y+7))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+50) && (lcd_pixel_x_address <= STEADY_X+57))&& (lcd_pixel_y_address == STEADY_Y+15))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
		   
						end
					/*End of Steady Screen for Game*/
					
					/*Bang Screen for Game*/
					else if (game_states == J_1_STATE || game_states == J_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		localparam BANG_X = 105;
		localparam BANG_Y = 150;
		localparam BANG_COLOUR = 16'h0000;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				if (((lcd_pixel_y_address >=BANG_Y+3) && (lcd_pixel_y_address <= BANG_Y+4))&& (lcd_pixel_x_address == BANG_X+7))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_y_address >=BANG_Y+10) && (lcd_pixel_y_address <= BANG_Y+12))&& (lcd_pixel_x_address == BANG_X+7))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y+7))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y+15))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+1))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+6))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+8))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+14))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+2))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+5))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+9))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+13))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				//Letter A
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+10))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=BANG_X+10) && (lcd_pixel_x_address <= BANG_X+17))&& (lcd_pixel_y_address == BANG_Y))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_x_address >=BANG_X+10) && (lcd_pixel_x_address <= BANG_X+17))&& (lcd_pixel_y_address == BANG_Y+7))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+17))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
					
				//Letter N
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+20))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+27))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+1))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+2))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+3))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
					
				
				else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+3))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+4))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+5))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+5))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+6))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+7))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end

				
				else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+7))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+8))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+9))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+9))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+10))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+11))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				
				
				else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+11))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+12))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+13))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				
				//Letter G
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+30))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=BANG_X+30) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_x_address >=BANG_X+34) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y+7))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_x_address >=BANG_X+30) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y+15))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_y_address >=BANG_Y+7) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+37))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end	
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
			
						end
					/*End of Bang Screen for Game*/
					
					/*Kill First Player for Game*/
					else if (game_states == L_1_STATE || game_states == L_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;


				if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+6)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+11)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+7)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+10)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
				//2P 
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
					
				
				else 	
					begin
						//lcd_pixel_data <= 16'hFFFF;
						lcd_pixel_data <= 16'hFFFF;
					end
			
						end
					/*End of Kill First Player for Game*/
					
					/*Kill Second Player for Game*/
					else if (game_states == K_1_STATE || game_states == K_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;


				if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
				//2P 
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+6)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+11)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+7)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+10)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				
				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
					
				
				else 	
					begin
						//lcd_pixel_data <= 16'hFFFF;
						lcd_pixel_data <= 16'hFFFF;
					end
				 
			
						end
					/*End of Kill Second Player for Game*/
					
					/*Kill Both Players for Game*/
					else if (game_states == M_1_STATE || game_states == M_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;


				if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+6)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+11)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+7)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+10)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
				//2P SELECTION SCREEN + 2nd Gunman
				
				//EXPLODE2d Head of GUNMAN2
				//GUNMAN2_X=100
				//GUNMAN2_Y=100
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+6)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+11)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+7)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+10)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				
				
				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
					
				
				else 	
					begin
						//lcd_pixel_data <= 16'hFFFF;
						lcd_pixel_data <= 16'hFFFF;
					end
				 
		   
						end
					/*End of Kill Both Players for Game*/
					
					/*First Player Winner for Game*/
					else if (game_states == Q_1_STATE || game_states == Q_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;


		localparam WINNER_X=80;
		localparam WINNER_Y=150;
		localparam WINNER_COLOUR=16'h0000;

		localparam _1P_X = 140;
		localparam _1P_Y = 150;
		localparam _1P_COLOUR = 16'h0000;

		/*
		localparam _2P_X = 140;
		localparam _2P_Y = 150;
		localparam _2P_COLOUR = 16'h0000;
		*/

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					

				
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+7))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//I	
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+14))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//N
				//Letter N
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+20))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+27))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+1))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+2))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+4))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+6))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end

				
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//N//Letter N
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+30))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+37))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+1))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+2))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+4))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+6))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end

				
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//E
				//Letter E
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+40))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y+7))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y+15))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//Letter R
				else if (((lcd_pixel_y_address >= WINNER_Y) && (lcd_pixel_y_address <= (WINNER_Y+15)))&& (lcd_pixel_x_address == WINNER_X+50))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=WINNER_X+50) && (lcd_pixel_x_address <= (WINNER_X+57)))&& (lcd_pixel_y_address == WINNER_Y))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= (WINNER_Y+7)))&& (lcd_pixel_x_address == (WINNER_X+57)))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= WINNER_X+50) && (lcd_pixel_x_address <= (WINNER_X+57)))&& (lcd_pixel_y_address == (WINNER_Y+7)))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+51) && (lcd_pixel_y_address==WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+52) && (lcd_pixel_y_address==WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+53) && (lcd_pixel_y_address==WINNER_Y+11)) 
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+54) && (lcd_pixel_y_address==WINNER_Y+12))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+55) && (lcd_pixel_y_address==WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+56) && (lcd_pixel_y_address==WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+57) && (lcd_pixel_y_address==WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end	
				
				//Player One
					//1
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+1))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+2))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+3))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==_1P_X+23) && (lcd_pixel_y_address == _1P_Y))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+23) && (lcd_pixel_y_address == _1P_Y+1))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+3))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+4))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+5))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
					
				else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= _1P_Y+15))&& (lcd_pixel_x_address == _1P_X+24))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=_1P_X+20) && (lcd_pixel_x_address <= _1P_X+28))&& (lcd_pixel_y_address == _1P_Y+15))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				//P	
				else if (((lcd_pixel_y_address >= _1P_Y) && (lcd_pixel_y_address <= (_1P_Y+15)))&& (lcd_pixel_x_address == _1P_X+10))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=_1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == _1P_Y))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= (_1P_Y+7)))&& (lcd_pixel_x_address == (_1P_X+17)))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= _1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == (_1P_Y+7)))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
					
				//PLAYER 2
			/*
				else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= _2P_Y+7))&& (lcd_pixel_x_address == _2P_X+27))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y+7))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y+15))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_y_address >=_2P_Y+8) && (lcd_pixel_y_address <= _2P_Y+15))&& (lcd_pixel_x_address == _2P_X+20))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >= _2P_Y) && (lcd_pixel_y_address <= (_2P_Y+15)))&& (lcd_pixel_x_address == _2P_X+10))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=_2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == _2P_Y))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= (_2P_Y+7)))&& (lcd_pixel_x_address == (_2P_X+17)))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= _2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == (_2P_Y+7)))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				//
				//
				*/
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
			
						end
					/*End of First Player Winner for Game*/
					
					/*Second Player Winner for Game*/
					else if (game_states == R_1_STATE || game_states == R_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;


		localparam WINNER_X=80;
		localparam WINNER_Y=150;
		localparam WINNER_COLOUR=16'h0000;

		localparam _2P_X = 140;
		localparam _2P_Y = 150;
		localparam _2P_COLOUR = 16'h0000;


		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					

				
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+7))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//I	
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+14))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//N
				//Letter N
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+20))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+27))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+1))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+2))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+4))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+6))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end

				
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//N//Letter N
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+30))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+37))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+1))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+2))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+4))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+6))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end

				
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//E
				//Letter E
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+40))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y+7))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y+15))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//Letter R
				else if (((lcd_pixel_y_address >= WINNER_Y) && (lcd_pixel_y_address <= (WINNER_Y+15)))&& (lcd_pixel_x_address == WINNER_X+50))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=WINNER_X+50) && (lcd_pixel_x_address <= (WINNER_X+57)))&& (lcd_pixel_y_address == WINNER_Y))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= (WINNER_Y+7)))&& (lcd_pixel_x_address == (WINNER_X+57)))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= WINNER_X+50) && (lcd_pixel_x_address <= (WINNER_X+57)))&& (lcd_pixel_y_address == (WINNER_Y+7)))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+51) && (lcd_pixel_y_address==WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+52) && (lcd_pixel_y_address==WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+53) && (lcd_pixel_y_address==WINNER_Y+11)) 
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+54) && (lcd_pixel_y_address==WINNER_Y+12))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+55) && (lcd_pixel_y_address==WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+56) && (lcd_pixel_y_address==WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+57) && (lcd_pixel_y_address==WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end	
				/*
				//Player One
					//1
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+1))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+2))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+3))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==_1P_X+23) && (lcd_pixel_y_address == _1P_Y))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+23) && (lcd_pixel_y_address == _1P_Y+1))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+3))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+4))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+5))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				
				else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= _1P_Y+15))&& (lcd_pixel_x_address == _1P_X+24))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=_1P_X+20) && (lcd_pixel_x_address <= _1P_X+28))&& (lcd_pixel_y_address == _1P_Y+15))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				//P	
				else if (((lcd_pixel_y_address >= _1P_Y) && (lcd_pixel_y_address <= (_1P_Y+15)))&& (lcd_pixel_x_address == _1P_X+10))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=_1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == _1P_Y))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= (_1P_Y+7)))&& (lcd_pixel_x_address == (_1P_X+17)))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= _1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == (_1P_Y+7)))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
				*/	
				
				
				//PLAYER 2
			
				else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= _2P_Y+7))&& (lcd_pixel_x_address == _2P_X+27))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y+7))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y+15))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_y_address >=_2P_Y+8) && (lcd_pixel_y_address <= _2P_Y+15))&& (lcd_pixel_x_address == _2P_X+20))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >= _2P_Y) && (lcd_pixel_y_address <= (_2P_Y+15)))&& (lcd_pixel_x_address == _2P_X+10))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=_2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == _2P_Y))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= (_2P_Y+7)))&& (lcd_pixel_x_address == (_2P_X+17)))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= _2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == (_2P_Y+7)))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				//
				//
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
		   
						end
					/*End of Second Player Winner for Game*/
					
					/*Next Screen for Player Two for Game*/
					else if (game_states == O_1_STATE || game_states == O_2_STATE)
						begin
							// LCD Display
							localparam LCD_WIDTH  = 240;
							localparam LCD_HEIGHT = 320;

							//1P
							localparam GUNMAN_X = 115;
							localparam GUNMAN_Y = 250;
							localparam BODY_COLOUR = 16'h0000;
							//localparam SCARF_COLOUR = 16'h07E0;
							localparam BELT_COLOUR = 16'hDA22;
							localparam GUN_COLOUR = 16'hA516;
							localparam PANTS_COLOUR = 16'h001F;
							localparam EXPLODE = 16'hF800;

							//2P
							localparam GUNMAN2_X = 115;
							localparam GUNMAN2_Y = 50;
							localparam BODY2_COLOUR = 16'h0000;
							//localparam SCARF2_COLOUR = 16'hF81F;
							localparam BELT2_COLOUR = 16'hDA22;
							localparam GUN2_COLOUR = 16'hA516;
							localparam PANTS2_COLOUR = 16'h001F;
							localparam EXPLODE2 = 16'hF800;

							localparam NEXT_X = 105;
							localparam NEXT_Y = 150;
							localparam NEXT_COLOUR = 16'h0000;
							
							if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+6)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+11)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+7)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+10)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							
							//Gunman Body
							
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end	
							
								
							//2P 
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
								
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							
							//GUNMAN2 Body
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end			
							
							//Letter N
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end

							
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							//Letter E
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+10))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+15))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							
							
							//Letter X
							//else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y-1))
							//	begin			
							//		lcd_pixel_data[15:0] <= NEXT_COLOUR;
							//	end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								

							
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end



							
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
								
							//else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y-1))
								//begin			
									//lcd_pixel_data[15:0] <= NEXT_COLOUR;
								//end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end		
								
							//Letter T
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+34))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+30) && (lcd_pixel_x_address <= NEXT_X+38))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else 	
								begin	
									lcd_pixel_data <= 16'hFFFF;
								end
					
						end
					/*End of Next Screen for Player Two for Game*/
					
					/*Next Screen for Player One for Game*/
					else if (game_states == N_1_STATE || game_states == N_2_STATE)
						begin
							// LCD Display
							//
							localparam LCD_WIDTH  = 240;
							localparam LCD_HEIGHT = 320;

							//1P
							localparam GUNMAN_X = 115;
							localparam GUNMAN_Y = 250;
							localparam BODY_COLOUR = 16'h0000;
							//localparam SCARF_COLOUR = 16'h07E0;
							localparam BELT_COLOUR = 16'hDA22;
							localparam GUN_COLOUR = 16'hA516;
							localparam PANTS_COLOUR = 16'h001F;
							localparam EXPLODE = 16'hF800;

							//2P
							localparam GUNMAN2_X = 115;
							localparam GUNMAN2_Y = 50;
							localparam BODY2_COLOUR = 16'h0000;
							//localparam SCARF2_COLOUR = 16'hF81F;
							localparam BELT2_COLOUR = 16'hDA22;
							localparam GUN2_COLOUR = 16'hA516;
							localparam PANTS2_COLOUR = 16'h001F;
							localparam EXPLODE2 = 16'hF800;

							localparam NEXT_X = 105;
							localparam NEXT_Y = 150;
							localparam NEXT_COLOUR = 16'h0000;
							
										//HEAD
							if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end

							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							
							//Gunman Body
							
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end	
							
								
							//2P 
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+6)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+11)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+7)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+10)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							
							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							
							//GUNMAN2 Body
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							//Letter N
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end

							
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							//Letter E
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+10))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+15))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							
							
							//Letter X
							//else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y-1))
							//	begin			
							//		lcd_pixel_data[15:0] <= NEXT_COLOUR;
							//	end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								

							
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end



							
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
								
							//else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y-1))
								//begin			
									//lcd_pixel_data[15:0] <= NEXT_COLOUR;
								//end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end		
								
							//Letter T
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+34))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+30) && (lcd_pixel_x_address <= NEXT_X+38))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else 	
								begin	
									lcd_pixel_data <= 16'hFFFF;
								end
							
						end
					/*End of Next Screen for Player One for Game*/
					
					/*Next Screen for Both Players for Game*/
					else if (game_states == P_1_STATE || game_states == P_2_STATE)
						begin
							// LCD Display
							//
							localparam LCD_WIDTH  = 240;
							localparam LCD_HEIGHT = 320;

							//1P
							localparam GUNMAN_X = 115;
							localparam GUNMAN_Y = 250;
							localparam BODY_COLOUR = 16'h0000;
							//localparam SCARF_COLOUR = 16'h07E0;
							localparam BELT_COLOUR = 16'hDA22;
							localparam GUN_COLOUR = 16'hA516;
							localparam PANTS_COLOUR = 16'h001F;
							localparam EXPLODE = 16'hF800;

							//2P
							localparam GUNMAN2_X = 115;
							localparam GUNMAN2_Y = 50;
							localparam BODY2_COLOUR = 16'h0000;
							//localparam SCARF2_COLOUR = 16'hF81F;
							localparam BELT2_COLOUR = 16'hDA22;
							localparam GUN2_COLOUR = 16'hA516;
							localparam PANTS2_COLOUR = 16'h001F;
							localparam EXPLODE2 = 16'hF800;

							localparam NEXT_X = 105;
							localparam NEXT_Y = 150;
							localparam NEXT_COLOUR = 16'h0000;
							
							if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+6)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+11)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+7)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+10)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							
							//Gunman Body
							
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end	
							
								
							//2P SELECTION SCREEN + 2nd Gunman
							
							//EXPLODE2d Head of GUNMAN2
							//GUNMAN2_X=100
							//GUNMAN2_Y=100
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+6)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+11)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+7)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+10)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							
							
							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							
							//GUNMAN2 Body
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end	
							//Letter N
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end

							
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							//Letter E
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+10))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+15))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							
							
							//Letter X
							//else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y-1))
							//	begin			
							//		lcd_pixel_data[15:0] <= NEXT_COLOUR;
							//	end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								

							
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end



							
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
								
							//else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y-1))
								//begin			
									//lcd_pixel_data[15:0] <= NEXT_COLOUR;
								//end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end		
								
							//Letter T
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+34))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+30) && (lcd_pixel_x_address <= NEXT_X+38))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							else 	
								begin	
									lcd_pixel_data <= 16'hFFFF;
								end
						
						end
					/*End of Next Screen for Both Players for Game*/
					
				end
				/* Player 1 ends. */
			
			else if ( PLAYER_ID == 2 )
				begin
					localparam SCARF2_COLOUR = 16'h07E0;
					localparam SCARF_COLOUR = 16'hF81F;
					
					/* Beginning of Main screen of the game. */
					if ( game_states == A_STATE  )
						begin
						
							localparam READY_X = 100;
							localparam READY_Y = 130;
							localparam READY_COLOUR = 16'hFFFF;
							localparam STEADY_X = 95;
							localparam STEADY_Y = 150;
							localparam STEADY_COLOUR = 16'hFFFF;
							localparam BANG_X = 105;
							localparam BANG_Y = 170;
							localparam BANG_COLOUR = 16'hFFFF;

							//1P
							localparam GUNMAN_X = 85;
							localparam GUNMAN_Y = 200;
							localparam BODY_COLOUR = 16'hFFFF;
							localparam BOX_COLOUR = 16'hFFFF;
							////localparam SCARF_COLOUR = 16'h07E0;
							localparam BELT_COLOUR = 16'hDA22;
							localparam GUN_COLOUR = 16'hA516;
							localparam PANTS_COLOUR = 16'h001F;
							localparam EXPLODE = 16'hF800;

							//2P
							localparam GUNMAN2_X = 145;
							localparam GUNMAN2_Y = 200;
							localparam BODY2_COLOUR = 16'hFFFF;
							localparam BOX2_COLOUR = 16'hFFFF;
							//localparam SCARF2_COLOUR = 16'hF81F;
							localparam BELT2_COLOUR = 16'hDA22;
							localparam GUN2_COLOUR = 16'hA516;
							localparam PANTS2_COLOUR = 16'h001F;
							localparam EXPLODE2 = 16'hF800;
							
							//WORD READY
							//READY=30
							
							//Letter R
							if (((lcd_pixel_y_address >= READY_Y) && (lcd_pixel_y_address <= (READY_Y+15)))&& (lcd_pixel_x_address == READY_X))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
								
							else if (((lcd_pixel_x_address >=READY_X) && (lcd_pixel_x_address <= (READY_X+7)))&& (lcd_pixel_y_address == READY_Y))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= (READY_Y+7)))&& (lcd_pixel_x_address == (READY_X+7)))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >= READY_X) && (lcd_pixel_x_address <= (READY_X+7)))&& (lcd_pixel_y_address == (READY_Y+7)))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if ((lcd_pixel_x_address==READY_X+1) && (lcd_pixel_y_address==READY_Y+9))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==READY_X+2) && (lcd_pixel_y_address==READY_Y+10))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==READY_X+3) && (lcd_pixel_y_address==READY_Y+11)) 
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==READY_X+4) && (lcd_pixel_y_address==READY_Y+12))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==READY_X+5) && (lcd_pixel_y_address==READY_Y+13))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==READY_X+6) && (lcd_pixel_y_address==READY_Y+14))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==READY_X+7) && (lcd_pixel_y_address==READY_Y+15))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	 
								end
								
							//Letter E
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+10))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y+7))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y+15))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
								
							//Letter A
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+20))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=READY_X+20) && (lcd_pixel_x_address <= READY_X+27))&& (lcd_pixel_y_address == READY_Y))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+20) && (lcd_pixel_x_address <= READY_X+27))&& (lcd_pixel_y_address == READY_Y+7))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+27))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
								
							//Letter D
							else if (((lcd_pixel_y_address >=READY_Y+4) && (lcd_pixel_y_address <= READY_Y+11))&& (lcd_pixel_x_address == READY_X+37))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+30))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+30) && (lcd_pixel_x_address <= READY_X+33))&& (lcd_pixel_y_address == READY_Y))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+30) && (lcd_pixel_x_address <= READY_X+33))&& (lcd_pixel_y_address == READY_Y+15))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if ((lcd_pixel_x_address==READY_X+33)  && (lcd_pixel_y_address==READY_Y))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if ((lcd_pixel_x_address==READY_X+33)  && (lcd_pixel_y_address==READY_Y+15))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if ((lcd_pixel_x_address==READY_X+34) && (lcd_pixel_y_address==READY_Y+1))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==READY_X+34) && (lcd_pixel_y_address==READY_Y+14))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==READY_X+35) && (lcd_pixel_y_address==READY_Y+2))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if ((lcd_pixel_x_address==READY_X+35) && (lcd_pixel_y_address==READY_Y+13))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if ((lcd_pixel_x_address==READY_X+36) && (lcd_pixel_y_address==READY_Y+3))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if ((lcd_pixel_x_address==READY_X+36) && (lcd_pixel_y_address==READY_Y+12))
								begin			
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							
							//Letter Y
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+47))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end	
							else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+7))&& (lcd_pixel_x_address == READY_X+40))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
								
							else if (((lcd_pixel_x_address >=READY_X+40) && (lcd_pixel_x_address <= READY_X+47))&& (lcd_pixel_y_address == READY_Y+7))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=READY_X+40) && (lcd_pixel_x_address <= READY_X+47))&& (lcd_pixel_y_address == READY_Y+15))
								begin
									lcd_pixel_data[15:0] <= READY_COLOUR;
								end
							
							
							//STEADY_Y+ & STEADY_X+
							//STEADY_COLOUR
							//Letter S
							//else
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+7))&& (lcd_pixel_x_address == STEADY_X))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y+7))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y+15))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=STEADY_Y+8) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+7))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
								
								//Letter T
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+14))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STEADY_X+10) && (lcd_pixel_x_address <= STEADY_X+17))&& (lcd_pixel_y_address == STEADY_Y))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							
							//Letter E
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+20))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y+7))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y+15))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							
							//Letter A
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+30))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STEADY_X+30) && (lcd_pixel_x_address <= STEADY_X+37))&& (lcd_pixel_y_address == STEADY_Y))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+30) && (lcd_pixel_x_address <= STEADY_X+37))&& (lcd_pixel_y_address == STEADY_Y+7))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+37))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
								
							//Letter D
							else if (((lcd_pixel_y_address >=STEADY_Y+4) && (lcd_pixel_y_address <= STEADY_Y+11))&& (lcd_pixel_x_address == STEADY_X+47))
								begin
									lcd_pixel_data[15:0] <=STEADY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+40))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+40) && (lcd_pixel_x_address <= STEADY_X+43))&& (lcd_pixel_y_address == STEADY_Y))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+40) && (lcd_pixel_x_address <= STEADY_X+43))&& (lcd_pixel_y_address == STEADY_Y+15))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+43) && (lcd_pixel_y_address == STEADY_Y))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==STEADY_X+43) && (lcd_pixel_y_address == STEADY_Y+15))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;	
								end
							else if ((lcd_pixel_x_address==STEADY_X+44) && (lcd_pixel_y_address == STEADY_Y+1))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+44) && (lcd_pixel_y_address == STEADY_Y+14))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+45) && (lcd_pixel_y_address == STEADY_Y+2))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+45) && (lcd_pixel_y_address == STEADY_Y+13))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+46) && (lcd_pixel_y_address == STEADY_Y+3))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if ((lcd_pixel_x_address==STEADY_X+46) && (lcd_pixel_y_address == STEADY_Y+12))
								begin			
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							
							//Letter Y
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+57))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end	
							else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+7))&& (lcd_pixel_x_address == STEADY_X+50))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
								
							else if (((lcd_pixel_x_address >=STEADY_X+50) && (lcd_pixel_x_address <= STEADY_X+57))&& (lcd_pixel_y_address == STEADY_Y+7))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STEADY_X+50) && (lcd_pixel_x_address <= STEADY_X+57))&& (lcd_pixel_y_address == STEADY_Y+15))
								begin
									lcd_pixel_data[15:0] <= STEADY_COLOUR;
								end
								
							
							//BANG_Y+=70
							//BANG_X+=30
							//BANG_COLOUR
							//Letter B
							else if (((lcd_pixel_y_address >=BANG_Y+3) && (lcd_pixel_y_address <= BANG_Y+4))&& (lcd_pixel_x_address == BANG_X+7))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_y_address >=BANG_Y+10) && (lcd_pixel_y_address <= BANG_Y+12))&& (lcd_pixel_x_address == BANG_X+7))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
								
							else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y+7))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y+15))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+1))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+6))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+8))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+14))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
								
							else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+2))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+5))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+9))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+13))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							//Letter A
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+10))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=BANG_X+10) && (lcd_pixel_x_address <= BANG_X+17))&& (lcd_pixel_y_address == BANG_Y))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_x_address >=BANG_X+10) && (lcd_pixel_x_address <= BANG_X+17))&& (lcd_pixel_y_address == BANG_Y+7))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+17))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
								
							//Letter N
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+20))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+27))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+1))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+2))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+3))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+3))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+4))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+5))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+5))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+6))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+7))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end

							
							else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+7))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+8))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+9))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+9))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+10))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+11))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							
							
							else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+11))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+12))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+13))
								begin			
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							
							
							//Letter G
							else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+30))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=BANG_X+30) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_x_address >=BANG_X+34) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y+7))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_x_address >=BANG_X+30) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y+15))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end
							else if (((lcd_pixel_y_address >=BANG_Y+7) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+37))
								begin
									lcd_pixel_data[15:0] <= BANG_COLOUR;
								end						
							
							//HEAD
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							
							//Gunman Body
							
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end	
								
							//HEAD
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							
							//GUNMAN2 Body
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end	
							else 	
								begin
									lcd_pixel_data <= 16'h0000;
								end
							
						end 
						/* End of Main screen of the game. */
					
					/*Selecting 1-Player Mode*/
					else if ( game_states == B_STATE )
						begin
						
						localparam LCD_WIDTH  = 240;
						localparam LCD_HEIGHT = 320;

						//1P
						localparam GUNMAN_X = 50;
						localparam GUNMAN_Y = 150;
						localparam BODY_COLOUR = 16'h0000;
						//localparam SCARF_COLOUR = 16'h07E0;
						localparam BELT_COLOUR = 16'hDA22;
						localparam GUN_COLOUR = 16'hA516;
						localparam PANTS_COLOUR = 16'h001F;
						localparam EXPLODE = 16'hF800;

						//2P
						localparam GUNMAN2_X = 130;
						localparam GUNMAN2_Y = 150;
						localparam BODY2_COLOUR = 16'h0000;
						//localparam SCARF2_COLOUR = 16'hF81F;
						localparam BELT2_COLOUR = 16'hDA22;
						localparam GUN2_COLOUR = 16'hA516;
						localparam PANTS2_COLOUR = 16'h001F;
						localparam EXPLODE2 = 16'hF800;


						localparam _1P_X = 53;
						localparam _1P_Y = 120;
						localparam _1P_COLOUR = 16'h0000;

						localparam _2P_X = 150;
						localparam _2P_Y = 120;
						localparam _2P_COLOUR = 16'h0000;

						localparam BOX_COLOUR = 16'h0000;
						localparam BOX2_COLOUR = 16'h0000;


								//Player One
									//1
								if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+1))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+2))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+3))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if ((lcd_pixel_x_address==_1P_X+3) && (lcd_pixel_y_address == _1P_Y))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+3) && (lcd_pixel_y_address == _1P_Y+1))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+3))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+4))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+5))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
									
								else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= _1P_Y+15))&& (lcd_pixel_x_address == _1P_X+4))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >=_1P_X) && (lcd_pixel_x_address <= _1P_X+8))&& (lcd_pixel_y_address == _1P_Y+15))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								//P	
								else if (((lcd_pixel_y_address >= _1P_Y) && (lcd_pixel_y_address <= (_1P_Y+15)))&& (lcd_pixel_x_address == _1P_X+10))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if (((lcd_pixel_x_address >=_1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == _1P_Y))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= (_1P_Y+7)))&& (lcd_pixel_x_address == (_1P_X+17)))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >= _1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == (_1P_Y+7)))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
									
								//PLAYER 2
							
								else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= _2P_Y+7))&& (lcd_pixel_x_address == _2P_X+7))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y+7))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y+15))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_y_address >=_2P_Y+8) && (lcd_pixel_y_address <= _2P_Y+15))&& (lcd_pixel_x_address == _2P_X))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_y_address >= _2P_Y) && (lcd_pixel_y_address <= (_2P_Y+15)))&& (lcd_pixel_x_address == _2P_X+10))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
									
								else if (((lcd_pixel_x_address >=_2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == _2P_Y))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= (_2P_Y+7)))&& (lcd_pixel_x_address == (_2P_X+17)))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >= _2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == (_2P_Y+7)))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								//
								//
								
								//Gunman 1
								
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end

								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT_COLOUR;
									end
								
								//Gunman Body
								
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end	
								
								//BOX for P1
								else if (((lcd_pixel_y_address >=(GUNMAN_Y-5)) && (lcd_pixel_y_address <= (GUNMAN_Y+38)))&&(lcd_pixel_x_address == (GUNMAN_X-8)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end	
								else if (((lcd_pixel_y_address >=(GUNMAN_Y-5)) && (lcd_pixel_y_address <= (GUNMAN_Y+38)))&&(lcd_pixel_x_address == (GUNMAN_X+26)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X-8) && (lcd_pixel_x_address <= (GUNMAN_X+26)))&&(lcd_pixel_y_address == (GUNMAN_Y-5)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X-8) && (lcd_pixel_x_address <= (GUNMAN_X+26)))&&(lcd_pixel_y_address == (GUNMAN_Y+38)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end	
									
								//2P 
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
							
								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								
								//GUNMAN2 Body
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end	
									
								//DUPLICATE FOR SELECTING OPTION	
										
								
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+47)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+50)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+47)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+50)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+45)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+52)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+45)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+52)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+48)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+49)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+46) && (lcd_pixel_x_address <= (GUNMAN2_X+51)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+46) && (lcd_pixel_x_address <= (GUNMAN2_X+51)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+48) && (lcd_pixel_x_address <= (GUNMAN2_X+49)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+48) && (lcd_pixel_x_address <= (GUNMAN2_X+49)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								
								//GUNMAN2 Body
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN2_X+39) && (lcd_pixel_x_address >= (GUNMAN2_X+38)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN2_X+39) && (lcd_pixel_x_address >= (GUNMAN2_X+38)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+58) && (lcd_pixel_x_address <= (GUNMAN2_X+59)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+58) && (lcd_pixel_x_address <= (GUNMAN2_X+59)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+37)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+36)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+60)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+61)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+40)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+41)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+42)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+43)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+56)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+57)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+54)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+44)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+45)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+52)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+53)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+42)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+43)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+41)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+54)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end	

								else 	
									begin
										//lcd_pixel_data <= 16'hFFFF;
										lcd_pixel_data <= 16'hFFFF;
									end

						end
					/*End of Selecting 1-Player Mode*/
					
					/*Selecting 2-Player Mode*/
					else if ( game_states == C_STATE )
						begin
											
						localparam LCD_WIDTH  = 240;
						localparam LCD_HEIGHT = 320;

						//1P
						localparam GUNMAN_X = 50;
						localparam GUNMAN_Y = 150;
						localparam BODY_COLOUR = 16'h0000;
						//localparam SCARF_COLOUR = 16'h07E0;
						localparam BELT_COLOUR = 16'hDA22;
						localparam GUN_COLOUR = 16'hA516;
						localparam PANTS_COLOUR = 16'h001F;
						localparam EXPLODE = 16'hF800;

						//2P
						localparam GUNMAN2_X = 130;
						localparam GUNMAN2_Y = 150;
						localparam BODY2_COLOUR = 16'h0000;
						//localparam SCARF2_COLOUR = 16'hF81F;
						localparam BELT2_COLOUR = 16'hDA22;
						localparam GUN2_COLOUR = 16'hA516;
						localparam PANTS2_COLOUR = 16'h001F;
						localparam EXPLODE2 = 16'hF800;


						localparam _1P_X = 53;
						localparam _1P_Y = 120;
						localparam _1P_COLOUR = 16'h0000;

						localparam _2P_X = 150;
						localparam _2P_Y = 120;
						localparam _2P_COLOUR = 16'h0000;

						localparam BOX_COLOUR = 16'h0000;
						localparam BOX2_COLOUR = 16'h0000;



								if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+1))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+2))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+2) && (lcd_pixel_y_address == _1P_Y+3))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if ((lcd_pixel_x_address==_1P_X+3) && (lcd_pixel_y_address == _1P_Y))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+3) && (lcd_pixel_y_address == _1P_Y+1))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+3))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+4))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								else if ((lcd_pixel_x_address==_1P_X+1) && (lcd_pixel_y_address == _1P_Y+5))
									begin			
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
									
								else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= _1P_Y+15))&& (lcd_pixel_x_address == _1P_X+4))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >=_1P_X) && (lcd_pixel_x_address <= _1P_X+8))&& (lcd_pixel_y_address == _1P_Y+15))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								//P	
								else if (((lcd_pixel_y_address >= _1P_Y) && (lcd_pixel_y_address <= (_1P_Y+15)))&& (lcd_pixel_x_address == _1P_X+10))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
									
								else if (((lcd_pixel_x_address >=_1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == _1P_Y))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= (_1P_Y+7)))&& (lcd_pixel_x_address == (_1P_X+17)))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >= _1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == (_1P_Y+7)))
									begin
										lcd_pixel_data[15:0] <= _1P_COLOUR;
									end	
									
								//PLAYER 2
							
								else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= _2P_Y+7))&& (lcd_pixel_x_address == _2P_X+7))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y+7))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_x_address >=_2P_X) && (lcd_pixel_x_address <= _2P_X+7))&& (lcd_pixel_y_address == _2P_Y+15))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_y_address >=_2P_Y+8) && (lcd_pixel_y_address <= _2P_Y+15))&& (lcd_pixel_x_address == _2P_X))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								else if (((lcd_pixel_y_address >= _2P_Y) && (lcd_pixel_y_address <= (_2P_Y+15)))&& (lcd_pixel_x_address == _2P_X+10))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
									
								else if (((lcd_pixel_x_address >=_2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == _2P_Y))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= (_2P_Y+7)))&& (lcd_pixel_x_address == (_2P_X+17)))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								else if (((lcd_pixel_x_address >= _2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == (_2P_Y+7)))
									begin
										lcd_pixel_data[15:0] <= _2P_COLOUR;
									end	
								//
								//
								
								//Gunman 1
								
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end

								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT_COLOUR;
									end
								
								//Gunman Body
								
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
									begin
										lcd_pixel_data[15:0] <= BODY_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= GUN_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS_COLOUR;
									end	
								
								/*//BOX for P1
								else if (((lcd_pixel_y_address >=(GUNMAN_Y-5)) && (lcd_pixel_y_address <= (GUNMAN_Y+38)))&&(lcd_pixel_x_address == (GUNMAN_X-8)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end	
								else if (((lcd_pixel_y_address >=(GUNMAN_Y-5)) && (lcd_pixel_y_address <= (GUNMAN_Y+38)))&&(lcd_pixel_x_address == (GUNMAN_X+26)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X-8) && (lcd_pixel_x_address <= (GUNMAN_X+26)))&&(lcd_pixel_y_address == (GUNMAN_Y-5)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN_X-8) && (lcd_pixel_x_address <= (GUNMAN_X+26)))&&(lcd_pixel_y_address == (GUNMAN_Y+38)))
									begin
										lcd_pixel_data[15:0] <= BOX_COLOUR;
									end*/	
									
								//2P 
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
							
								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								
								//GUNMAN2 Body
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end	
									
								//DUPLICATE FOR SELECTING OPTION	
										
								
								//HEAD
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+47)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+50)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+47)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+50)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+45)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+52)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+44)) && (lcd_pixel_x_address <= (GUNMAN2_X+45)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=(GUNMAN2_X+52)) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+48)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+49)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								//green scarf h07E0
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+46) && (lcd_pixel_x_address <= (GUNMAN2_X+51)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+46) && (lcd_pixel_x_address <= (GUNMAN2_X+51)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+48) && (lcd_pixel_x_address <= (GUNMAN2_X+49)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+48) && (lcd_pixel_x_address <= (GUNMAN2_X+49)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= SCARF2_COLOUR;
									end	
									
								//brown belt
								//DA22
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BELT2_COLOUR;
									end
								
								//GUNMAN2 Body
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+40) && (lcd_pixel_x_address <= (GUNMAN2_X+57)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+44) && (lcd_pixel_x_address <= (GUNMAN2_X+53)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
									
								//Arms
								else if (((lcd_pixel_x_address <=GUNMAN2_X+39) && (lcd_pixel_x_address >= (GUNMAN2_X+38)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address <=GUNMAN2_X+39) && (lcd_pixel_x_address >= (GUNMAN2_X+38)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_x_address >=GUNMAN2_X+58) && (lcd_pixel_x_address <= (GUNMAN2_X+59)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X+58) && (lcd_pixel_x_address <= (GUNMAN2_X+59)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end	
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+37)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+36)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+60)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+61)))
									begin
										lcd_pixel_data[15:0] <= BODY2_COLOUR;
									end
								
								
								
								//silver guns
								//A516
								//left
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+40)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+41)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+42)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+43)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								//right
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+56)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+57)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+54)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= GUN2_COLOUR;
									end
									
								//blue legs h001F
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+44)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+45)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+52)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+53)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
									
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+42)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+43)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+41)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+54)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+55)))
									begin
										lcd_pixel_data[15:0] <= PANTS2_COLOUR;
									end	
								
								//BOX for P2
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y-5)) && (lcd_pixel_y_address <= (GUNMAN2_Y+38)))&&(lcd_pixel_x_address == (GUNMAN2_X-8)))
									begin
										lcd_pixel_data[15:0] <= BOX2_COLOUR;
									end	
								else if (((lcd_pixel_y_address >=(GUNMAN2_Y-5)) && (lcd_pixel_y_address <= (GUNMAN2_Y+38)))&&(lcd_pixel_x_address == (GUNMAN2_X+66)))
									begin
										lcd_pixel_data[15:0] <= BOX2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X-8) && (lcd_pixel_x_address <= (GUNMAN2_X+66)))&&(lcd_pixel_y_address == (GUNMAN2_Y-5)))
									begin
										lcd_pixel_data[15:0] <= BOX2_COLOUR;
									end
								else if (((lcd_pixel_x_address >=GUNMAN2_X-8) && (lcd_pixel_x_address <= (GUNMAN2_X+66)))&&(lcd_pixel_y_address == (GUNMAN2_Y+38)))
									begin
										lcd_pixel_data[15:0] <= BOX2_COLOUR;
									end
									
								
								else 	
									begin
										//lcd_pixel_data <= 16'hFFFF;
										lcd_pixel_data <= 16'hFFFF;
									end
								  
							
											
									
						end
					/*End of Selecting 2-Player Mode*/
					
					/* Beginning of Select Player screen. */
					else if ( game_states == D_1_STATE || game_states == D_2_STATE  )
						begin
						
							localparam LCD_WIDTH  = 240;
							localparam LCD_HEIGHT = 320;

							localparam STARTGAME_X = 105;
							localparam STARTGAME_Y = 150;
							localparam STARTGAME_COLOUR = 16'h0000;

							//1P
							localparam GUNMAN_X = 115;
							localparam GUNMAN_Y = 250;
							localparam BODY_COLOUR = 16'h0000;
							//localparam SCARF_COLOUR = 16'h07E0;
							localparam BELT_COLOUR = 16'hDA22;
							localparam GUN_COLOUR = 16'hA516;
							localparam PANTS_COLOUR = 16'h001F;
							localparam EXPLODE = 16'hF800;

							//2P
							localparam GUNMAN2_X = 115;
							localparam GUNMAN2_Y = 50;
							localparam BODY2_COLOUR = 16'h0000;
							//localparam SCARF2_COLOUR = 16'hF81F;
							localparam BELT2_COLOUR = 16'hDA22;
							localparam GUN2_COLOUR = 16'hA516;
							localparam PANTS2_COLOUR = 16'h001F;
							localparam EXPLODE2 = 16'hF800;
							
							//STARTGAME_Y+ & STARTGAME_X+
							//STARTGAME_COLOUR
							//Letter S
							//else
							if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= STARTGAME_Y+7))&& (lcd_pixel_x_address == STARTGAME_X))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STARTGAME_X) && (lcd_pixel_x_address <= STARTGAME_X+7))&& (lcd_pixel_y_address == STARTGAME_Y))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STARTGAME_X) && (lcd_pixel_x_address <= STARTGAME_X+7))&& (lcd_pixel_y_address == STARTGAME_Y+7))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STARTGAME_X) && (lcd_pixel_x_address <= STARTGAME_X+7))&& (lcd_pixel_y_address == STARTGAME_Y+15))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if (((lcd_pixel_y_address >=STARTGAME_Y+8) && (lcd_pixel_y_address <= STARTGAME_Y+15))&& (lcd_pixel_x_address == STARTGAME_X+7))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
								
								//Letter T
							else if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= STARTGAME_Y+15))&& (lcd_pixel_x_address == STARTGAME_X+14))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STARTGAME_X+10) && (lcd_pixel_x_address <= STARTGAME_X+17))&& (lcd_pixel_y_address == STARTGAME_Y))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							
							
							//Letter A
							else if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= STARTGAME_Y+15))&& (lcd_pixel_x_address == STARTGAME_X+20))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STARTGAME_X+20) && (lcd_pixel_x_address <= STARTGAME_X+27))&& (lcd_pixel_y_address == STARTGAME_Y))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if (((lcd_pixel_x_address >=STARTGAME_X+20) && (lcd_pixel_x_address <= STARTGAME_X+27))&& (lcd_pixel_y_address == STARTGAME_Y+7))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= STARTGAME_Y+15))&& (lcd_pixel_x_address == STARTGAME_X+27))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
								
							//Letter R
							else if (((lcd_pixel_y_address >= STARTGAME_Y) && (lcd_pixel_y_address <= (STARTGAME_Y+15)))&& (lcd_pixel_x_address == STARTGAME_X+30))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
								
							else if (((lcd_pixel_x_address >=STARTGAME_X+30) && (lcd_pixel_x_address <= (STARTGAME_X+37)))&& (lcd_pixel_y_address == STARTGAME_Y))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= (STARTGAME_Y+7)))&& (lcd_pixel_x_address == (STARTGAME_X+37)))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end	
							else if (((lcd_pixel_x_address >= STARTGAME_X+30) && (lcd_pixel_x_address <= (STARTGAME_X+37)))&& (lcd_pixel_y_address == (STARTGAME_Y+7)))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+31) && (lcd_pixel_y_address==STARTGAME_Y+9))
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+32) && (lcd_pixel_y_address==STARTGAME_Y+10))
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+33) && (lcd_pixel_y_address==STARTGAME_Y+11)) 
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+34) && (lcd_pixel_y_address==STARTGAME_Y+12))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+35) && (lcd_pixel_y_address==STARTGAME_Y+13))
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+36) && (lcd_pixel_y_address==STARTGAME_Y+14))
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	 
								end
							else if ((lcd_pixel_x_address==STARTGAME_X+37) && (lcd_pixel_y_address==STARTGAME_Y+15))
								begin			
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;	 
								end
							//Letter T
							else if (((lcd_pixel_y_address >=STARTGAME_Y) && (lcd_pixel_y_address <= STARTGAME_Y+15))&& (lcd_pixel_x_address == STARTGAME_X+44))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=STARTGAME_X+40) && (lcd_pixel_x_address <= STARTGAME_X+47))&& (lcd_pixel_y_address == STARTGAME_Y))
								begin
									lcd_pixel_data[15:0] <= STARTGAME_COLOUR;
								end
							
							
							//HEAD
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end

							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							
							//Gunman Body
							
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end	
							
								
								
							
							//HEAD
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//scarf 
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							
							//GUNMAN2 Body
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end	
							else 	
								begin	
									lcd_pixel_data <= 16'hFFFF;
								end
							
						end 
						/* End of Select Player screen. */
					
					/*In-Between Screens*/
					else if ( game_states == E_1_STATE || game_states == G_1_STATE || game_states == I_1_STATE || game_states == E_2_STATE || game_states == G_2_STATE || game_states == I_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				//HEAD
				if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
		   
						
						end
					/*End of In-Between Screens*/
					
					/*Ready Screen for Game*/
					else if ( game_states == F_1_STATE || game_states == F_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		localparam READY_X = 105;
		localparam READY_Y = 150;
		localparam READY_COLOUR = 16'h0000;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				//Letter R
				if (((lcd_pixel_y_address >= READY_Y) && (lcd_pixel_y_address <= (READY_Y+15)))&& (lcd_pixel_x_address == READY_X))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=READY_X) && (lcd_pixel_x_address <= (READY_X+7)))&& (lcd_pixel_y_address == READY_Y))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= (READY_Y+7)))&& (lcd_pixel_x_address == (READY_X+7)))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= READY_X) && (lcd_pixel_x_address <= (READY_X+7)))&& (lcd_pixel_y_address == (READY_Y+7)))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if ((lcd_pixel_x_address==READY_X+1) && (lcd_pixel_y_address==READY_Y+9))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==READY_X+2) && (lcd_pixel_y_address==READY_Y+10))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==READY_X+3) && (lcd_pixel_y_address==READY_Y+11)) 
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==READY_X+4) && (lcd_pixel_y_address==READY_Y+12))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==READY_X+5) && (lcd_pixel_y_address==READY_Y+13))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==READY_X+6) && (lcd_pixel_y_address==READY_Y+14))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==READY_X+7) && (lcd_pixel_y_address==READY_Y+15))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	 
					end
					
				//Letter E
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+10))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y+7))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+10) && (lcd_pixel_x_address <= READY_X+17))&& (lcd_pixel_y_address == READY_Y+15))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
					
				//Letter A
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+20))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=READY_X+20) && (lcd_pixel_x_address <= READY_X+27))&& (lcd_pixel_y_address == READY_Y))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+20) && (lcd_pixel_x_address <= READY_X+27))&& (lcd_pixel_y_address == READY_Y+7))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+27))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
					
				//Letter D
				else if (((lcd_pixel_y_address >=READY_Y+4) && (lcd_pixel_y_address <= READY_Y+11))&& (lcd_pixel_x_address == READY_X+37))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+30))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+30) && (lcd_pixel_x_address <= READY_X+33))&& (lcd_pixel_y_address == READY_Y))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+30) && (lcd_pixel_x_address <= READY_X+33))&& (lcd_pixel_y_address == READY_Y+15))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if ((lcd_pixel_x_address==READY_X+33)  && (lcd_pixel_y_address==READY_Y))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if ((lcd_pixel_x_address==READY_X+33)  && (lcd_pixel_y_address==READY_Y+15))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if ((lcd_pixel_x_address==READY_X+34) && (lcd_pixel_y_address==READY_Y+1))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==READY_X+34) && (lcd_pixel_y_address==READY_Y+14))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==READY_X+35) && (lcd_pixel_y_address==READY_Y+2))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if ((lcd_pixel_x_address==READY_X+35) && (lcd_pixel_y_address==READY_Y+13))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if ((lcd_pixel_x_address==READY_X+36) && (lcd_pixel_y_address==READY_Y+3))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if ((lcd_pixel_x_address==READY_X+36) && (lcd_pixel_y_address==READY_Y+12))
					begin			
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				
				//Letter Y
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+15))&& (lcd_pixel_x_address == READY_X+47))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end	
				else if (((lcd_pixel_y_address >=READY_Y) && (lcd_pixel_y_address <= READY_Y+7))&& (lcd_pixel_x_address == READY_X+40))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=READY_X+40) && (lcd_pixel_x_address <= READY_X+47))&& (lcd_pixel_y_address == READY_Y+7))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=READY_X+40) && (lcd_pixel_x_address <= READY_X+47))&& (lcd_pixel_y_address == READY_Y+15))
					begin
						lcd_pixel_data[15:0] <= READY_COLOUR;
					end
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
			
						end
					/*End of Ready Screen for Game*/
					
					/*Steady Screen for Game*/
					else if (game_states == H_1_STATE || game_states == H_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		localparam STEADY_X = 105;
		localparam STEADY_Y = 150;
		localparam STEADY_COLOUR = 16'h0000;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+7))&& (lcd_pixel_x_address == STEADY_X))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y+7))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X) && (lcd_pixel_x_address <= STEADY_X+7))&& (lcd_pixel_y_address == STEADY_Y+15))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=STEADY_Y+8) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+7))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
					
					//Letter T
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+14))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=STEADY_X+10) && (lcd_pixel_x_address <= STEADY_X+17))&& (lcd_pixel_y_address == STEADY_Y))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				
				//Letter E
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+20))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y+7))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+20) && (lcd_pixel_x_address <= STEADY_X+27))&& (lcd_pixel_y_address == STEADY_Y+15))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				
				//Letter A
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+30))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=STEADY_X+30) && (lcd_pixel_x_address <= STEADY_X+37))&& (lcd_pixel_y_address == STEADY_Y))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+30) && (lcd_pixel_x_address <= STEADY_X+37))&& (lcd_pixel_y_address == STEADY_Y+7))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+37))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
					
				//Letter D
				else if (((lcd_pixel_y_address >=STEADY_Y+4) && (lcd_pixel_y_address <= STEADY_Y+11))&& (lcd_pixel_x_address == STEADY_X+47))
					begin
						lcd_pixel_data[15:0] <=STEADY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+40))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+40) && (lcd_pixel_x_address <= STEADY_X+43))&& (lcd_pixel_y_address == STEADY_Y))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+40) && (lcd_pixel_x_address <= STEADY_X+43))&& (lcd_pixel_y_address == STEADY_Y+15))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+43) && (lcd_pixel_y_address == STEADY_Y))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==STEADY_X+43) && (lcd_pixel_y_address == STEADY_Y+15))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;	
					end
				else if ((lcd_pixel_x_address==STEADY_X+44) && (lcd_pixel_y_address == STEADY_Y+1))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+44) && (lcd_pixel_y_address == STEADY_Y+14))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+45) && (lcd_pixel_y_address == STEADY_Y+2))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+45) && (lcd_pixel_y_address == STEADY_Y+13))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+46) && (lcd_pixel_y_address == STEADY_Y+3))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if ((lcd_pixel_x_address==STEADY_X+46) && (lcd_pixel_y_address == STEADY_Y+12))
					begin			
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				
				//Letter Y
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+15))&& (lcd_pixel_x_address == STEADY_X+57))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end	
				else if (((lcd_pixel_y_address >=STEADY_Y) && (lcd_pixel_y_address <= STEADY_Y+7))&& (lcd_pixel_x_address == STEADY_X+50))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=STEADY_X+50) && (lcd_pixel_x_address <= STEADY_X+57))&& (lcd_pixel_y_address == STEADY_Y+7))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=STEADY_X+50) && (lcd_pixel_x_address <= STEADY_X+57))&& (lcd_pixel_y_address == STEADY_Y+15))
					begin
						lcd_pixel_data[15:0] <= STEADY_COLOUR;
					end
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
		   
						end
					/*End of Steady Screen for Game*/
					
					/*Bang Screen for Game*/
					else if (game_states == J_1_STATE || game_states == J_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		localparam BANG_X = 105;
		localparam BANG_Y = 150;
		localparam BANG_COLOUR = 16'h0000;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				if (((lcd_pixel_y_address >=BANG_Y+3) && (lcd_pixel_y_address <= BANG_Y+4))&& (lcd_pixel_x_address == BANG_X+7))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_y_address >=BANG_Y+10) && (lcd_pixel_y_address <= BANG_Y+12))&& (lcd_pixel_x_address == BANG_X+7))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y+7))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_x_address >=BANG_X) && (lcd_pixel_x_address <= BANG_X+4))&& (lcd_pixel_y_address == BANG_Y+15))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+1))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+6))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+8))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+5) && (lcd_pixel_y_address == BANG_Y+14))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+2))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+5))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+9))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+6) && (lcd_pixel_y_address == BANG_Y+13))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				//Letter A
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+10))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=BANG_X+10) && (lcd_pixel_x_address <= BANG_X+17))&& (lcd_pixel_y_address == BANG_Y))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_x_address >=BANG_X+10) && (lcd_pixel_x_address <= BANG_X+17))&& (lcd_pixel_y_address == BANG_Y+7))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+17))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
					
				//Letter N
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+20))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+27))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+1))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+2))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+21) && (lcd_pixel_y_address == BANG_Y+3))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
					
				
				else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+3))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+4))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+22) && (lcd_pixel_y_address == BANG_Y+5))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+5))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+6))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+23) && (lcd_pixel_y_address == BANG_Y+7))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end

				
				else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+7))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+8))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+24) && (lcd_pixel_y_address == BANG_Y+9))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+9))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+10))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+25) && (lcd_pixel_y_address == BANG_Y+11))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				
				
				else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+11))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+12))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if ((lcd_pixel_x_address==BANG_X+26) && (lcd_pixel_y_address == BANG_Y+13))
					begin			
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				
				
				//Letter G
				else if (((lcd_pixel_y_address >=BANG_Y) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+30))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=BANG_X+30) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_x_address >=BANG_X+34) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y+7))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_x_address >=BANG_X+30) && (lcd_pixel_x_address <= BANG_X+37))&& (lcd_pixel_y_address == BANG_Y+15))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end
				else if (((lcd_pixel_y_address >=BANG_Y+7) && (lcd_pixel_y_address <= BANG_Y+15))&& (lcd_pixel_x_address == BANG_X+37))
					begin
						lcd_pixel_data[15:0] <= BANG_COLOUR;
					end	
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
			
						end
					/*End of Bang Screen for Game*/
					
					/*Kill First Player for Game*/
					else if (game_states == L_1_STATE || game_states == L_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;


				if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+6)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+11)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+7)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+10)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
				//2P 
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
					
				
				else 	
					begin
						//lcd_pixel_data <= 16'hFFFF;
						lcd_pixel_data <= 16'hFFFF;
					end
			
						end
					/*End of Kill First Player for Game*/
					
					/*Kill Second Player for Game*/
					else if (game_states == K_1_STATE || game_states == K_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;


				if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
				//2P 
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+6)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+11)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+7)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+10)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				
				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
					
				
				else 	
					begin
						//lcd_pixel_data <= 16'hFFFF;
						lcd_pixel_data <= 16'hFFFF;
					end
				 
			
						end
					/*End of Kill Second Player for Game*/
					
					/*Kill Both Players for Game*/
					else if (game_states == M_1_STATE || game_states == M_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;


				if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+6)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+11)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+7)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+10)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE;
					end
				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
				//2P SELECTION SCREEN + 2nd Gunman
				
				//EXPLODE2d Head of GUNMAN2
				//GUNMAN2_X=100
				//GUNMAN2_Y=100
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+6)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+11)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+7)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+10)))
					begin
						lcd_pixel_data[15:0] <= EXPLODE2;
					end
				
				
				
				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
					
				
				else 	
					begin
						//lcd_pixel_data <= 16'hFFFF;
						lcd_pixel_data <= 16'hFFFF;
					end
				 
		   
						end
					/*End of Kill Both Players for Game*/
					
					/*First Player Winner for Game*/
					else if (game_states == Q_1_STATE || game_states == Q_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;


		localparam WINNER_X=80;
		localparam WINNER_Y=150;
		localparam WINNER_COLOUR=16'h0000;

		localparam _1P_X = 140;
		localparam _1P_Y = 150;
		localparam _1P_COLOUR = 16'h0000;

		/*
		localparam _2P_X = 140;
		localparam _2P_Y = 150;
		localparam _2P_COLOUR = 16'h0000;
		*/

		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					

				
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+7))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//I	
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+14))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//N
				//Letter N
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+20))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+27))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+1))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+2))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+4))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+6))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end

				
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//N//Letter N
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+30))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+37))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+1))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+2))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+4))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+6))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end

				
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//E
				//Letter E
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+40))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y+7))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y+15))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//Letter R
				else if (((lcd_pixel_y_address >= WINNER_Y) && (lcd_pixel_y_address <= (WINNER_Y+15)))&& (lcd_pixel_x_address == WINNER_X+50))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=WINNER_X+50) && (lcd_pixel_x_address <= (WINNER_X+57)))&& (lcd_pixel_y_address == WINNER_Y))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= (WINNER_Y+7)))&& (lcd_pixel_x_address == (WINNER_X+57)))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= WINNER_X+50) && (lcd_pixel_x_address <= (WINNER_X+57)))&& (lcd_pixel_y_address == (WINNER_Y+7)))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+51) && (lcd_pixel_y_address==WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+52) && (lcd_pixel_y_address==WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+53) && (lcd_pixel_y_address==WINNER_Y+11)) 
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+54) && (lcd_pixel_y_address==WINNER_Y+12))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+55) && (lcd_pixel_y_address==WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+56) && (lcd_pixel_y_address==WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+57) && (lcd_pixel_y_address==WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end	
				
				//Player One
					//1
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+1))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+2))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+3))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==_1P_X+23) && (lcd_pixel_y_address == _1P_Y))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+23) && (lcd_pixel_y_address == _1P_Y+1))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+3))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+4))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+5))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
					
				else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= _1P_Y+15))&& (lcd_pixel_x_address == _1P_X+24))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=_1P_X+20) && (lcd_pixel_x_address <= _1P_X+28))&& (lcd_pixel_y_address == _1P_Y+15))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				//P	
				else if (((lcd_pixel_y_address >= _1P_Y) && (lcd_pixel_y_address <= (_1P_Y+15)))&& (lcd_pixel_x_address == _1P_X+10))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=_1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == _1P_Y))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= (_1P_Y+7)))&& (lcd_pixel_x_address == (_1P_X+17)))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= _1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == (_1P_Y+7)))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
					
				//PLAYER 2
			/*
				else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= _2P_Y+7))&& (lcd_pixel_x_address == _2P_X+27))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y+7))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y+15))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_y_address >=_2P_Y+8) && (lcd_pixel_y_address <= _2P_Y+15))&& (lcd_pixel_x_address == _2P_X+20))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >= _2P_Y) && (lcd_pixel_y_address <= (_2P_Y+15)))&& (lcd_pixel_x_address == _2P_X+10))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=_2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == _2P_Y))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= (_2P_Y+7)))&& (lcd_pixel_x_address == (_2P_X+17)))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= _2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == (_2P_Y+7)))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				//
				//
				*/
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
			
						end
					/*End of First Player Winner for Game*/
					
					/*Second Player Winner for Game*/
					else if (game_states == R_1_STATE || game_states == R_2_STATE)
						begin
						
		localparam LCD_WIDTH  = 240;
		localparam LCD_HEIGHT = 320;


		localparam WINNER_X=80;
		localparam WINNER_Y=150;
		localparam WINNER_COLOUR=16'h0000;

		localparam _2P_X = 140;
		localparam _2P_Y = 150;
		localparam _2P_COLOUR = 16'h0000;


		//1P
		localparam GUNMAN_X = 115;
		localparam GUNMAN_Y = 250;
		localparam BODY_COLOUR = 16'h0000;
		//localparam SCARF_COLOUR = 16'h07E0;
		localparam BELT_COLOUR = 16'hDA22;
		localparam GUN_COLOUR = 16'hA516;
		localparam PANTS_COLOUR = 16'h001F;
		localparam EXPLODE = 16'hF800;

		//2P
		localparam GUNMAN2_X = 115;
		localparam GUNMAN2_Y = 50;
		localparam BODY2_COLOUR = 16'h0000;
		//localparam SCARF2_COLOUR = 16'hF81F;
		localparam BELT2_COLOUR = 16'hDA22;
		localparam GUN2_COLOUR = 16'hA516;
		localparam PANTS2_COLOUR = 16'h001F;
		localparam EXPLODE2 = 16'hF800;

				if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X) && (lcd_pixel_y_address == WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+1) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+2) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+3) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					

				
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+4) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+5) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+6) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+7) && (lcd_pixel_y_address == WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+7))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//I	
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+14))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//N
				//Letter N
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+20))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+27))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+1))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+2))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+21) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+4))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+22) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+6))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+23) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end

				
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+24) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+25) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+26) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//N//Letter N
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+30))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+37))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+1))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+2))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+31) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+3))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+4))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+32) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+5))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+6))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+33) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end

				
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+7))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+8))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+34) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+35) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				
				
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+11))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+12))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+36) && (lcd_pixel_y_address == WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//E
				//Letter E
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= WINNER_Y+15))&& (lcd_pixel_x_address == WINNER_X+40))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y+7))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if (((lcd_pixel_x_address >=WINNER_X+40) && (lcd_pixel_x_address <= WINNER_X+47))&& (lcd_pixel_y_address == WINNER_Y+15))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				//Letter R
				else if (((lcd_pixel_y_address >= WINNER_Y) && (lcd_pixel_y_address <= (WINNER_Y+15)))&& (lcd_pixel_x_address == WINNER_X+50))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=WINNER_X+50) && (lcd_pixel_x_address <= (WINNER_X+57)))&& (lcd_pixel_y_address == WINNER_Y))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=WINNER_Y) && (lcd_pixel_y_address <= (WINNER_Y+7)))&& (lcd_pixel_x_address == (WINNER_X+57)))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= WINNER_X+50) && (lcd_pixel_x_address <= (WINNER_X+57)))&& (lcd_pixel_y_address == (WINNER_Y+7)))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;
					end
				else if ((lcd_pixel_x_address==WINNER_X+51) && (lcd_pixel_y_address==WINNER_Y+9))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+52) && (lcd_pixel_y_address==WINNER_Y+10))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+53) && (lcd_pixel_y_address==WINNER_Y+11)) 
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+54) && (lcd_pixel_y_address==WINNER_Y+12))
					begin
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+55) && (lcd_pixel_y_address==WINNER_Y+13))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	
					end
				else if ((lcd_pixel_x_address==WINNER_X+56) && (lcd_pixel_y_address==WINNER_Y+14))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end
				else if ((lcd_pixel_x_address==WINNER_X+57) && (lcd_pixel_y_address==WINNER_Y+15))
					begin			
						lcd_pixel_data[15:0] <= WINNER_COLOUR;	 
					end	
				/*
				//Player One
					//1
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+1))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+2))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+22) && (lcd_pixel_y_address == _1P_Y+3))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==_1P_X+23) && (lcd_pixel_y_address == _1P_Y))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+23) && (lcd_pixel_y_address == _1P_Y+1))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+3))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+4))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				else if ((lcd_pixel_x_address==_1P_X+21) && (lcd_pixel_y_address == _1P_Y+5))
					begin			
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				
				else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= _1P_Y+15))&& (lcd_pixel_x_address == _1P_X+24))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=_1P_X+20) && (lcd_pixel_x_address <= _1P_X+28))&& (lcd_pixel_y_address == _1P_Y+15))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				//P	
				else if (((lcd_pixel_y_address >= _1P_Y) && (lcd_pixel_y_address <= (_1P_Y+15)))&& (lcd_pixel_x_address == _1P_X+10))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=_1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == _1P_Y))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=_1P_Y) && (lcd_pixel_y_address <= (_1P_Y+7)))&& (lcd_pixel_x_address == (_1P_X+17)))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= _1P_X+10) && (lcd_pixel_x_address <= (_1P_X+17)))&& (lcd_pixel_y_address == (_1P_Y+7)))
					begin
						lcd_pixel_data[15:0] <= _1P_COLOUR;
					end	
				*/	
				
				
				//PLAYER 2
			
				else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= _2P_Y+7))&& (lcd_pixel_x_address == _2P_X+27))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y+7))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_x_address >=_2P_X+20) && (lcd_pixel_x_address <= _2P_X+27))&& (lcd_pixel_y_address == _2P_Y+15))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				else if (((lcd_pixel_y_address >=_2P_Y+8) && (lcd_pixel_y_address <= _2P_Y+15))&& (lcd_pixel_x_address == _2P_X+20))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >= _2P_Y) && (lcd_pixel_y_address <= (_2P_Y+15)))&& (lcd_pixel_x_address == _2P_X+10))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
					
				else if (((lcd_pixel_x_address >=_2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == _2P_Y))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=_2P_Y) && (lcd_pixel_y_address <= (_2P_Y+7)))&& (lcd_pixel_x_address == (_2P_X+17)))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				else if (((lcd_pixel_x_address >= _2P_X+10) && (lcd_pixel_x_address <= (_2P_X+17)))&& (lcd_pixel_y_address == (_2P_Y+7)))
					begin
						lcd_pixel_data[15:0] <= _2P_COLOUR;
					end	
				//
				//
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end

				
				//green scarf h07E0
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT_COLOUR;
					end
				
				//Gunman Body
				
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS_COLOUR;
					end	
				
					
					
				
				//HEAD
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//scarf 
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= SCARF2_COLOUR;
					end	
					
				//brown belt
				//DA22
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BELT2_COLOUR;
					end
				
				//GUNMAN2 Body
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
					
				//Arms
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end	
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
					begin
						lcd_pixel_data[15:0] <= BODY2_COLOUR;
					end
				
				
				
				//silver guns
				//A516
				//left
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				//right
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= GUN2_COLOUR;
					end
					
				//blue legs h001F
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
					
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end
				else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
					begin
						lcd_pixel_data[15:0] <= PANTS2_COLOUR;
					end	
				else 	
					begin	
						lcd_pixel_data <= 16'hFFFF;
					end
		   
						end
					/*End of Second Player Winner for Game*/
					
					/*Next Screen for Player Two for Game*/
					else if (game_states == O_1_STATE || game_states == O_2_STATE)
						begin
							// LCD Display
							localparam LCD_WIDTH  = 240;
							localparam LCD_HEIGHT = 320;

							//1P
							localparam GUNMAN_X = 115;
							localparam GUNMAN_Y = 250;
							localparam BODY_COLOUR = 16'h0000;
							//localparam SCARF_COLOUR = 16'h07E0;
							localparam BELT_COLOUR = 16'hDA22;
							localparam GUN_COLOUR = 16'hA516;
							localparam PANTS_COLOUR = 16'h001F;
							localparam EXPLODE = 16'hF800;

							//2P
							localparam GUNMAN2_X = 115;
							localparam GUNMAN2_Y = 50;
							localparam BODY2_COLOUR = 16'h0000;
							//localparam SCARF2_COLOUR = 16'hF81F;
							localparam BELT2_COLOUR = 16'hDA22;
							localparam GUN2_COLOUR = 16'hA516;
							localparam PANTS2_COLOUR = 16'h001F;
							localparam EXPLODE2 = 16'hF800;

							localparam NEXT_X = 105;
							localparam NEXT_Y = 150;
							localparam NEXT_COLOUR = 16'h0000;
							
							if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+6)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+11)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+7)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+10)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							
							//Gunman Body
							
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end	
							
								
							//2P 
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+6)))
								
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+7)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+10)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+4)) && (lcd_pixel_x_address <= (GUNMAN2_X+5)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN2_X+12)) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+8)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							
							//GUNMAN2 Body
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end			
							
							//Letter N
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end

							
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							//Letter E
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+10))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+15))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							
							
							//Letter X
							//else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y-1))
							//	begin			
							//		lcd_pixel_data[15:0] <= NEXT_COLOUR;
							//	end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								

							
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end



							
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
								
							//else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y-1))
								//begin			
									//lcd_pixel_data[15:0] <= NEXT_COLOUR;
								//end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end		
								
							//Letter T
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+34))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+30) && (lcd_pixel_x_address <= NEXT_X+38))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else 	
								begin	
									lcd_pixel_data <= 16'hFFFF;
								end
					
						end
					/*End of Next Screen for Player Two for Game*/
					
					/*Next Screen for Player One for Game*/
					else if (game_states == N_1_STATE || game_states == N_2_STATE)
						begin
							// LCD Display
							//
							localparam LCD_WIDTH  = 240;
							localparam LCD_HEIGHT = 320;

							//1P
							localparam GUNMAN_X = 115;
							localparam GUNMAN_Y = 250;
							localparam BODY_COLOUR = 16'h0000;
							//localparam SCARF_COLOUR = 16'h07E0;
							localparam BELT_COLOUR = 16'hDA22;
							localparam GUN_COLOUR = 16'hA516;
							localparam PANTS_COLOUR = 16'h001F;
							localparam EXPLODE = 16'hF800;

							//2P
							localparam GUNMAN2_X = 115;
							localparam GUNMAN2_Y = 50;
							localparam BODY2_COLOUR = 16'h0000;
							//localparam SCARF2_COLOUR = 16'hF81F;
							localparam BELT2_COLOUR = 16'hDA22;
							localparam GUN2_COLOUR = 16'hA516;
							localparam PANTS2_COLOUR = 16'h001F;
							localparam EXPLODE2 = 16'hF800;

							localparam NEXT_X = 105;
							localparam NEXT_Y = 150;
							localparam NEXT_COLOUR = 16'h0000;
							
										//HEAD
							if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+6)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+7)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+5)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+7)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+10)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+2)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+1)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+4)) && (lcd_pixel_x_address <= (GUNMAN_X+5)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=(GUNMAN_X+12)) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+8)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end

							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							
							//Gunman Body
							
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end	
							
								
							//2P 
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+6)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+11)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+7)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+10)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							
							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							
							//GUNMAN2 Body
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							//Letter N
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end

							
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							//Letter E
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+10))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+15))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							
							
							//Letter X
							//else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y-1))
							//	begin			
							//		lcd_pixel_data[15:0] <= NEXT_COLOUR;
							//	end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								

							
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end



							
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
								
							//else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y-1))
								//begin			
									//lcd_pixel_data[15:0] <= NEXT_COLOUR;
								//end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end		
								
							//Letter T
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+34))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+30) && (lcd_pixel_x_address <= NEXT_X+38))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else 	
								begin	
									lcd_pixel_data <= 16'hFFFF;
								end
							
						end
					/*End of Next Screen for Player One for Game*/
					
					/*Next Screen for Both Players for Game*/
					else if (game_states == P_1_STATE || game_states == P_2_STATE)
						begin
							// LCD Display
							//
							localparam LCD_WIDTH  = 240;
							localparam LCD_HEIGHT = 320;

							//1P
							localparam GUNMAN_X = 115;
							localparam GUNMAN_Y = 250;
							localparam BODY_COLOUR = 16'h0000;
							//localparam SCARF_COLOUR = 16'h07E0;
							localparam BELT_COLOUR = 16'hDA22;
							localparam GUN_COLOUR = 16'hA516;
							localparam PANTS_COLOUR = 16'h001F;
							localparam EXPLODE = 16'hF800;

							//2P
							localparam GUNMAN2_X = 115;
							localparam GUNMAN2_Y = 50;
							localparam BODY2_COLOUR = 16'h0000;
							//localparam SCARF2_COLOUR = 16'hF81F;
							localparam BELT2_COLOUR = 16'hDA22;
							localparam GUN2_COLOUR = 16'hA516;
							localparam PANTS2_COLOUR = 16'h001F;
							localparam EXPLODE2 = 16'hF800;

							localparam NEXT_X = 105;
							localparam NEXT_Y = 150;
							localparam NEXT_COLOUR = 16'h0000;
							
							if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+3)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+7)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+6)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+11)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y)) && (lcd_pixel_y_address <= (GUNMAN_Y+10)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+7)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+8)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+9)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+3)) && (lcd_pixel_y_address <= (GUNMAN_Y+7)))&&(lcd_pixel_x_address == (GUNMAN_X+10)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE;
								end
							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+6) && (lcd_pixel_x_address <= (GUNMAN_X+11)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+8) && (lcd_pixel_x_address <= (GUNMAN_X+9)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT_COLOUR;
								end
							
							//Gunman Body
							
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X) && (lcd_pixel_x_address <= (GUNMAN_X+17)))&&(lcd_pixel_y_address == (GUNMAN_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+4) && (lcd_pixel_x_address <= (GUNMAN_X+13)))&&(lcd_pixel_y_address == (GUNMAN_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN_X-1) && (lcd_pixel_x_address >= (GUNMAN_X-2)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN_X+18) && (lcd_pixel_x_address <= (GUNMAN_X+19)))&&(lcd_pixel_y_address == (GUNMAN_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+19)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+24)))&&(lcd_pixel_x_address == (GUNMAN_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+23)) && (lcd_pixel_y_address <= (GUNMAN_Y+28)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+25)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN_Y+32)) && (lcd_pixel_y_address <= (GUNMAN_Y+33)))&&(lcd_pixel_x_address == (GUNMAN_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS_COLOUR;
								end	
							
								
							//2P SELECTION SCREEN + 2nd Gunman
							
							//EXPLODE2d Head of GUNMAN2
							//GUNMAN2_X=100
							//GUNMAN2_Y=100
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+3)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+7)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+6)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+11)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y)) && (lcd_pixel_y_address <= (GUNMAN2_Y+10)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+7)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+8)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+9)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+3)) && (lcd_pixel_y_address <= (GUNMAN2_Y+7)))&&(lcd_pixel_x_address == (GUNMAN2_X+10)))
								begin
									lcd_pixel_data[15:0] <= EXPLODE2;
								end
							
							
							
							
							//green scarf h07E0
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+6) && (lcd_pixel_x_address <= (GUNMAN2_X+11)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+8) && (lcd_pixel_x_address <= (GUNMAN2_X+9)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= SCARF2_COLOUR;
								end	
								
							//brown belt
							//DA22
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BELT2_COLOUR;
								end
							
							//GUNMAN2 Body
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+14)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+15)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X) && (lcd_pixel_x_address <= (GUNMAN2_X+17)))&&(lcd_pixel_y_address == (GUNMAN2_Y+16)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+19)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+22)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+23)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+4) && (lcd_pixel_x_address <= (GUNMAN2_X+13)))&&(lcd_pixel_y_address == (GUNMAN2_Y+24)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
								
							//Arms
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address <=GUNMAN2_X-1) && (lcd_pixel_x_address >= (GUNMAN2_X-2)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+17)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_x_address >=GUNMAN2_X+18) && (lcd_pixel_x_address <= (GUNMAN2_X+19)))&&(lcd_pixel_y_address == (GUNMAN2_Y+18)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end	
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-3)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X-4)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+20)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+19)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+21)))
								begin
									lcd_pixel_data[15:0] <= BODY2_COLOUR;
								end
							
							
							
							//silver guns
							//A516
							//left
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+0)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							//right
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+16)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+24)))&&(lcd_pixel_x_address == (GUNMAN2_X+17)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+23)) && (lcd_pixel_y_address <= (GUNMAN2_Y+28)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= GUN2_COLOUR;
								end
								
							//blue legs h001F
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+4)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+5)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+12)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+25)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+13)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
								
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+2)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+3)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+1)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+14)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end
							else if (((lcd_pixel_y_address >=(GUNMAN2_Y+32)) && (lcd_pixel_y_address <= (GUNMAN2_Y+33)))&&(lcd_pixel_x_address == (GUNMAN2_X+15)))
								begin
									lcd_pixel_data[15:0] <= PANTS2_COLOUR;
								end	
							//Letter N
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+1) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+2) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+3) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end

							
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+4) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+5) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+6) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							//Letter E
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+10))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+7))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if (((lcd_pixel_x_address >=NEXT_X+10) && (lcd_pixel_x_address <= NEXT_X+17))&& (lcd_pixel_y_address == NEXT_Y+15))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							
							
							//Letter X
							//else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y-1))
							//	begin			
							//		lcd_pixel_data[15:0] <= NEXT_COLOUR;
							//	end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+20) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+21) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+22) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+6))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+23) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								

							
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+7))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+8))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+24) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+9))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+10))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+4))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+25) && (lcd_pixel_y_address == NEXT_Y+5))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							
							
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+11))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+12))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+2))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+26) && (lcd_pixel_y_address == NEXT_Y+3))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end



							
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+13))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+14))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+15))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
								
							//else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y-1))
								//begin			
									//lcd_pixel_data[15:0] <= NEXT_COLOUR;
								//end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
							else if ((lcd_pixel_x_address==NEXT_X+27) && (lcd_pixel_y_address == NEXT_Y+1))
								begin			
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end		
								
							//Letter T
							else if (((lcd_pixel_y_address >=NEXT_Y) && (lcd_pixel_y_address <= NEXT_Y+15))&& (lcd_pixel_x_address == NEXT_X+34))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end	
							else if (((lcd_pixel_x_address >=NEXT_X+30) && (lcd_pixel_x_address <= NEXT_X+38))&& (lcd_pixel_y_address == NEXT_Y))
								begin
									lcd_pixel_data[15:0] <= NEXT_COLOUR;
								end
								
							else 	
								begin	
									lcd_pixel_data <= 16'hFFFF;
								end
						
						end
					/*End of Next Screen for Both Players for Game*/
				end
				/* Player 2 ends. */
			
		end
			
endmodule																		// End of the module.



